XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��PpP��w|���)�UE&�݁����.V��u�t�T%���20�<M�Z�fH�]�$�FD��k�S,Mݱ�t��E�F^ݶ��b��s�r��u^�Y���p#���6}�c��|8;[�pVB/���)�mQ1�V���m��yq���W����kg_񵑓$���`��p͢��QL<ߋ�A�P��������+*2�E��ȼK��:��\��n[�8��S�TH��II}	�]Ai.ǉ����%VS
 �3��y^�{�A)��*	<�PG���l�L��{���T�E�MХ@�)�48|��r�P0}kZ`r3h���$��	r��Yb���rL<+4&'��6���Me��7I��I߽���A^��� C��e08�Cv?ə���N�j^7,6��%{T}��F���|9���{����RSP���
WT���3R���Zq�&� ��r��Ǹ#��z~9a���|��x��2��4`LQE'��?}��s�����y{pEu�� (Z��3��|vR��>øN�Hv�{��Z6�ą�p���G��W��آ��UhA�$���	Bv&c�Cm5�cQ�Z��E ��uh'�Q�i�'���lۍ_d���<�C���T�q��,��<������O��nS��n�l |���UHkW�����D0>�nG��F%G��Ĕa-_{I���'��W��bm�|�d�Zk��F���q�����z0HA��©�ؼT����d�!�:�-�ϥ$L��O�1XlxVHYEB    9de1    1670
�?n̊�>�����: ��+U�|�}BIVA���Ɋ2�3��VE��e+�yxI�*XKl(�>I�j��jU����.�(���A�J(�b�y��-�H�`��Ĭu����^�!�� ش�6��b�z���x�C����[�;��bO��w	M�D� !�*v����$K=���SȗB�P*��)P�Fɴ�]�!��7�!����5(1X.Hk9�K|@��+ KSH�,��\#8?����$����R����k*�m�C������_rh?G��qI�+y	}0�Yg@\,���)�k�u��I��ZgI/��YaS^0o��!��_�Up�}>��ͨ��e]��b�O*��J�_X�D]��Mh2G|�=L<�
����p$S��;��@���}Q�`Zo)���r���3�jƄ�k]6�o��(��Сbt��~�6���h�X5~����.�ܖ�i��%A_����n�����A��� ��7÷�ڕd�["x�w��ء
 :�7�F�935�ׅJ���`��xXv���aƸ�랾�T����ə�s��o,�?�K�I�Ub�N�l�4T�|Agk;K6��eA�{�4��\]?t�5��䏈ο4#� ���������\��js'����Q�i<D���V���|��nJ����f�5Cc q-�����G������J@��N[o�����Hf�*�N�����L�Wl8��X�����zF�7��ޒDĐ��v�j�R���2b[��P�
�@Ng� ���*��$��C&�'��F�B*�r���Y�"�HwM��2hd�|�ґ�Ԫ�h�� ����P�&n*�-b_A��R�H�7ۍ����4�be.)��"�'��g�g��7K�=�oP�v�H���w�M|��ǥ�7�&cJ���G�����(ŦSy�%��颥�{'9v�����σ�ˊ��=�^I����^f��|d�x���/��ٗ��ϡ���\6y�)| �v���d��9��"d�;�*����Apyefi��Q�=��}�X�����_j���m�T�.�f�#O>�.b����s=6���/4h��o"7�v��ڠ���ҧ����M��2��ٸ�O|^^�(���J*8@c����f��������]_gk<�܈J�L�ah�;�^�'B���[v�y�`�٘K���^�9�{71��f�NI�n�����nV%#���]�@��r����}��2���n��D8t7�d�`ALwR�S����d���7k�lmx����`8�A���:��
��n�Um�&'/ڕ1A�~�FY��\4@ُ֡���I���G�7�	r���"EO��)��6*_��;���ԛ�S�C�܀3� �����n����J46�_���6��l����^8 i������.��4��+�C.�������l �n-*�\��L�ڸ��:E@=�n�-�$���EFw�w?���Tzy�ws&�v��=�	m�1����+3餉O�?���3m�%/��#v2.��l+�I:������.ߜ��pf���-�)��?����������S��G`�n1B3�ds5���eS�}'���ڪ�9��D��S&��Z~�������X)���ēc5������kt�����`�୐�2$�-���`�y|�2��IWt��h��WwVN�Q-z�d��F �����t��^�1_�s��3@ε�7��`�96�Vbh,��޸w|=�0�;+?+>d~�W�5�����ᡖ�����&�\>�Z�� �PS��~��zv ��E�҂���VzH�+*>6(�j"Y�_a�V����yD�0h���מ ]D���q3v�֕���R�\l�G�\��)�o�I�3�sUv�"�v=���̿kP�%�g����f��`�؍8�	���,�0�#)�?q�_�Ţ���A/0R�ϗ���A��4��H�6��+�}��\{���"S��h�J�'��B�[�b箄�ʺm� )��?�s��0R������ʜ\�(	�E�#�������HJ��&R����LZ���f�yW��P�Ɔ-�Zw�)wL�Tw����d2ЁIi@I)G?�q��ßW�QGV~��<PO<�&�iW�7�ba�nC�c��g6�)�V�X��}2�:$�s�� 0N�"���.���2@ΩIy?����`
i��P�Ww��z��O��a~�@������:���(uDV�tc��%8eBYW�4���V������&?�i�M6uVQ���D�ϧ���`�2̳��W�^�s	\�~�X�v%Y5����u7�(��ܑa����Nzz.��������}�j�3�f�&,�.�'���1�"�}��.7=>*�6xZ�¦��ª\�b����L���'�u;���&QJ]�75�\]�4v����~*��e�B�no/�&��?ou�3����%��h��^�ڏJ��+�Y�xȣQ�~H��s�����RP�,��?��M]<�4�_��+�*��YN� Ne%%�A�/@�2h\�����X; v��u�#?-�Ǿ����� �"�K+n��<���lbp���U�&��y��i����~���������a\|�@�S��K�E���`���<�q�+�����ܚ���`*n�m.���ޑ�|��~������*+�7'3p��k���?)�V�=
ʴ���k8Ǫ� h�wV*C�C��d���p��߲�_#"evp.#aɕh�J1R7�4RUwTu"b�zH��A�a2f$�4D6@��Z���c���a��^���#< �FcoƝU&7	㛭2� ��)!���wD��f(���w���G2욜����k������N�
�<����_�}�f��.�M�E��.=�q����7��Tp��&�'��#)���^�s�5�U$��|��䥈��-l���" *�=M�/҄�ʝI�qA_����f� ��xe��<�36�] v�,l&�.�G�X �r��f_k��OO���`�I	��o�L��/�8vs��G�)mM�\���~��D�\�,�(��#����<�?u�V_��w�_�ν�B�c���H�#I/�ғ��q�,/��}�Z��YX���<�3��)7�����V^#�Yo���P�~� �y�����r�P�1u�6��`M�j��9Z��FY�I%�LJh��ܚ"�̿��8�|��t������*��MA�g��D#΄ԣ�p����&���)�] ԰�� @�,��`�smbF����z���V�"���u��
���;������,eA����K'۶d3�㭧v�8��~u6��C<��x,�I���ɇ��z����F_�YJ6���aTUޞ�
�T���G{k�Bܽ��|1Ա�V��������R�M�/[�m�������]��,�� ��T�3�34_J,�0�_�w�?��4"yP��  tX�Ƨ��v����ӈ ��ԨՂu9��@9�+2�c��4?�_!��5���� �q���ƂD&ފ���ؙ��1<��B��zk��x��V ��}q��NKjƬI�\��U�*�e°D��0>��J�����������	aq�l�4�J*��+�?7p�z�cW�������y��'�V&Q{��;��˞�'D�� �����H �w�]���GYR-�˓�v�ٱ�r���C�-}&�f��+���=�ổ?��6u,�3s��2�̩���4�J�	5��/�����S�(GC[W�.r/M:S�}�u
L=)q1�'�ۣq�j�l/���a���k�,p
"���^��WE�����,�D���&&�l2MO�s"ѓE�!i�«���V���T̟�Ќ�JQ�A�d�s}�XB���AAW��/�7�4�#ŋN㲸��s3�����ɢ�eɟ�v�,��3~$���&��P�\l>/���/�v������ �������4H��E�����1�ґh���� NO(j(ۃn����P����Ǿ���#��&ߊ��nSGND����o�cwʚD���J�Q�����!�����ʾֆ���!�ڈK�	;ڲB���S�;�4��fC6i��)9�>e�vR�ċBY�8m�$��l�D��\nb��tم.4��^*hnE�h?���Ih��l�@��&��n>kc�Y���@�()�}�*�L�t+�^o����+�M{8+���[�;��+�＄\�_]���P�u�t�g������Q��|���9NX;PHu����]��HKwטޞJU�s>
_:�1칯\� _R�i}�d��M�a4��d���9���yũ�T�!� �NB"o����6` R>��dtZ�w�<��8�^��F��r�,<�\��j� 1k�D���}_>��VLM!(H�_�wX'�J���
 gM��4�0V�������vJc=b����~#���}Y)����4�'�(	�<%:�/�B�� ��q���Q��5��)Y0���| �/�1������X*�՞����bhKI�
��	K���G���O��)cr���獰2�1.��U�TQ�������&�c��@�I�����%���<��O�ͷo<�f-8�-��:�d[�Y����Pŵ�6vy���:s��9�TwT�#��hf��YҨ=�~^�4d��u0�V�_��E��dW��]���C��?���(_4�i���I�j�7y�'������W)L��$��H����1�����$tKE.^�������)=�r��6EHi�wugB���`a��YI4ɴ��)i4H���1X�:!-H�Pw�گ}��	� h$M���] �e�Z�}�4vq���F��;б����`�)���
�E5C����Y�)Τ�	�$P{�HH��������p$X�L�9`�7���ޣ^�������r�|^��h��3�Q,�}��N"�f$xQ9)�&*橫��oj��(��*��	�S��V���� 5�>��XO��:<�H���d�9v2�l���@���5a�"V�}�H����+��4P����/��m1��TY��6���wӑk�]�rޮ?v���v�	��.��iLU)G�+^�N*6 ."�-

9�0c�i��!!:޸>���#3K��4���
�fВάK���L�u�!X�7OE���=��RQ���fL�K�[�_\cՕ���2`���϶��G�^�::��]� 2�u�O��ġ�EQ�����<�^�TN�3�V��~ϵ�����?W�g�?
L�8�6��;laz�y��)�RONm��k�x�`�u��M|�|�lv o�S[�$橆�~�-.�q��]������`P/!����p����f�,xC���&|�h��>�=nE�築˜��,Ԑ����	�*Tѵ�1}�@�1m���o'��00�£"�o������r���~�96"���E9�bv����O��8�w�b]���u��x�1eG�8f�ÜB2ư��s���*bz8���8��%�8t}P�(z���"��c\�������W�(O��-�:*&�vz�r�%'�����lS#�Ȱ���2~�י�tMaT�&t�Aӑ��������{@U�o�p�L]Oi���EI�r��#��Q	�^��8ܭ}:|�[{�9���O�w�D�ߎ�V�){�p��& ����(�rJu���l�����+