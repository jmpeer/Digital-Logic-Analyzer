XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ǅ�ơ�ˇ_0���㝒 �	�"��ö��Y��`|tv�?fZF�k�+��B,bA��T����Qn��ǫ��ח���r�m�³�tie�=gpB��P}F��j*S+ӉD��a��|@�Ƥ��^uo# _��`�0 ���
QM��)�����G���:���.�#���z,u�"͟��kM�(�:W"�v��̋�`�T��'#'A��[mMd"�Pڥ��o6�ܖ�yJ^vwqE�8��D�S�^`#B��G��z��.��n�>	~xu��y4�j�`En���ā\C���[��>����i���N�Z�Vs��";A�Y�kW���h�K��Ƃ�����3���wu�ԩK@����j�;��u{�m.��.��A���<�������=d<wMvU�����p@]S�r�������|������x3����\�&6�De�~wV�ta�ِ쎴�$È���( �Q�m�;�ݠ�مȿ��;�H��8aP�a�Gr�-��mҸ��7UɕHZs�ͤCC�TyT�'��m`�y@7&�܁�iTE����vN��8�@�0���7��p�
n"��'8����[~iiD�A|��0����/{����[k����t��UʹQQdt�-o���0��Me����p��8���a�2@�����Z���e�d�cCçH$��A�]��m�4
nL��%7��M�FK��ۋ��T���K���Zõ�S�HQ��
H��[��M��oj��(7��4h<%}z����w'ר�ی�xXlxVHYEB    fa00    1f80>���ʻ�i����-l�L͘���	JJ� �
@B9~���.�euw�	ZYn�q"����NSz���Zt������8fCM�Kc��/ݸwmg�\����_Jc���z����=PVS�����A��񥇈�����܁��͆�j="*����9��G�E�k�c�?j�O{��-�E�vLIj�'l�`	�ӌ1���0�0 �M�WqP ��g��z����̧Zy����q�Ӡ��<��4���+q���$5�.������q\C���[6��h�	0�\,B��s@��_ 6`�z��\a۲X�$rɥ�>��E���Trh��	������(HR('���/3����~�8k �IW�>e,� xy�Ux�sl��g�la}[�	P;K��-���T��gO�薁�nɀ�;d��t.Gl�V�f����u-"�_����F'�V��fFn�V9[���˖R%.�C����T��&#),W�U^���~cd��t8-�>�� G�?�k��ݠd��&���@J�� #5-O���<���i�
����GU6��${�_J�>^��,��"Z���}�V��f���I�{e��%��r����Va6�"ɨ͑�ȣ�����2��mK�5��1�}���Y��ȭ�
��?^��}M��ආo�'tC��l�,���_��0���"�����V����p���=����« N�ǌ��f��cl0\�a[�ެvE_\�o	*��x��ۧ���M�!k����Jo�����2�Lޙ��p3g�`'�����\˾x'�rƻ4}�p��d���D�b�:AL�]�n������n��)�����TcЪ�3/��Pgjm�¢�i9�|V�ܣZN��rS�r�,"h��>����9���'@8P��q0geY*Ʒ��/C"�è��j�u��]aSg�kZ�'�Aڸ�؉5�X^'�X�G'�����"����y��fK
�%�@�ؕ0~>�44_Cfm�8����H�s�\�`9�2%�Cߠ?~�M,�˫o^��j���u	{������lrFl�4����m���]�^!	�s�߁�B~��1��Y�:��u�Q�Kvh�6�h�\�m/	-���=\��iy=0.����U��HrЙ�Q\�'h1�MG����"�]5���O��;񇥥�{����p �v����c\�!~��Q�&����҉q�0z���N]h?2H1�vܽ ����H�4>Rf�u��u�����:n2k�Ilw�2F�Ȥ``��tO�m^����U�C'q���isP鬲�ױ�؇&�_�pOvQ��U2�h����ׁ��o���J���
�x��	z�7��	0���`��7]4�ËͲ�q�[�F��Iv>���N[N���|_�R"����Nڛ�ѭ�Mm.��r
����`�L��(!��D�O��8���V��"M���Z��=�*8��o7JV�M�U4�+#۷�e7R��tdu$x��������&�~c,�u]3}~��i��LG0}g���*uw5�`�?.؜@�0K��RUOc��DȬ%�$z���\.P����W��\�q�u����ڱ		�i��"1����<�"6�m��������y���nr���ͪ4U<F;,�{��&��c�N���'�R�6�{V��Oz����tc��d����O�۱� v�:����ǔ �
J�h������k$���M��'7�2F�&�O���j�H�Oc>����A������jΓdIܬ���S�br�,Ҿ(���F��Ŀ�r�8�p�D��[A�n׸���k��#a/�;�;w��8��4#�
�:㇉-B1i��^i˞���<�>�k�ީ�K]����{5�(���N��8��*�i�Ut"�H�!��U5!��B�o������ 
J�#�j�ρO"K�88�"ޓ�8h�>�F�oW�?�����nv^a��-4i�"9�A[�&j�YHUB�3���ԉixK̏<i3Rߛ�#�����pz��h�v��j���dAF�v�����K�=����j�g0«����A"q��q�����ʷ�E<�Y�z��ϗ��Rfͥۥ*�ĭ�h�f�"����hh��w�)��l���F�?��p����Qv-K|�_��'�	44���?y���چ��G��uN����S?s��Q4�N;��e�q�A-KU���>�KH�O�|�]Mȫ����� W���IN%�ybH��=ռW?�^ǹ��e�hivJ����Sp��QL���n;�G��#B�}F�$�'fخ(N�>����RE6��l�+���^qd~�J4��ӭ���Q���_#,o!�퓑��IL�>�s˸.#���x�����.�� u����}wa��^"��FB���x�5������b����;޼)D)��y�b���X��\W:P�I�>쳞�zu��	���ƍH�ֆq/�*]+�V��VI���.�;^ /7�?֧� ��J�eq�k�3P*�d��&wn�uSɔ���k���e<,�osᏉ,�eP�s?y2,�f6�";�?��:?�H���@.`�O�)�ב��)��ܝ���J���|�����9��D�e�c%+��-��ǋ�s����@2�x�%o� q���G�����I['��턽�>�����uK���h_���q�jB+_s�Vj�@��~M��,H.~�lEq��`&���%/veV�O�Mmr�	���\t�;؉� ���,�d�}��U�j$�$�v��ǃ|�#m�F�1�À�lHO�/#��Jt{���L�v�L��&��T��ME�D~K#���KO���s�[卮���*A[�RH�S�/G���I����0ݺ������"���=�]=)�DΈ ?~�l[��h�oP^YU>E��Gv��w����X��u������=��LT?2�資��^�� �	��uC��^�D9�4��R�h��M`��gڝZ�D-�8��V	n��pE�M�A�*E;Uw!I�_�E4[;��-2�k�,��Kӷ޺n�b��-;RկR�8$V�-� 8�VPq�h���νҴ�	ȓ�Q�(�	,0 ��D>jƱ/[�����w� =���B��������c�=i�A��W�lo�F\q�+�������QF*/�h��Ԝ�T�Z_!�0��1ܲ	��@��"\ k$�ɸ�1ƠħK���c��0�@Cxd�7��`j�i0d	��f�eW�sN�����P��J���K���n� ��Qz�,��*I�pS�n���"���+�W�Ώ�$�0�\�C\7u�N7����|���;e�o$���Qq�T���+\2��KJ']8n��e��h�Ƚ�!��d��m�l���)��</�~�������e2��^m��/)߀�`�����`�qD@��B�?:��-�vZ�esme<4;ú���s�-@��~>]�T�7Y��g`M.aPR�"1���泙ʸ��#��ӀO{3Kg{�ɰ�3cx��?�Ȝ0\��c�|�8��/D�o����G�w���<�|�C�k��ub�	�a��W�C_���@.1�3XF���w��ߕ�7р��W D�8�"D��f89�4�����HVT�?�})<�5\�Vؖ^-ܗD7���i��8ͫ^�77�ǟ��d�H��ǻ���n��'~�<̹� ��)|Q��A�ƝJ�z�31p.Ǩ��Ნv�͌��`�ȡry�g���6��"LI�`�����IR�ӑ��f�|�k���:�FP3,FҊp9�#b�ȍ����
M��L"�l-�,��Ф�F��
9��&���b�y�X�0�	$@��05�2U���N���/���~���+���$�La|I���c�(6�+׆����u�t��(0���LE��Fl9ٕ�+�&�?w����4`��_�����\�h��'�B9�~:�k�8���@�?��Q)�F�:I�!*�2�+����-j8#�^Be+Q�\�� $�%rO�Ro�����lZ�u���Z��}@����r��D�<��6�(��/�#q�o�,��"�"0���r<�{����`����MzbZ��({"�`W"��/\��>�s��Y!�MHg��%�G�7�oI�L�������˕����$a��5��n�����Ym�'��^tF_���ՄE����&�{�A�''`Wu;��*8\�B���G�KZ���,�	��	�g��-��~=s)q�UQ�M�P����ĨAל�L���-F� ��j#��L���n��`��Hχ�؛�ՙ����i}v�WCO�'�G������x�)K�N��K&���G�r�ʁb��"�!9�6{�;��Ѭq�ʷ~��,k���Fᇹ�a�~�,���0}���BVM�*�|���� �?7YU)� ��c��*�-v�+Sr�xF���Δ��r�0��0����?<�7>�>���.�Pq�i��p/ĩzO�G�
L����ð5Y�@D�����dJ�ַ�}���,�n؁J���Rx&>��
g�����K/X�c�d:���d�9i8����z�o�;=�ZB1.��V�>��֌���m������nbǠ�L�����a��# J|,��gµ#�F�b��J�6c�P�2
	�5Jn�b+���7b�5)>���]T<e:����R�7�4-!apz��HnD@H��z�ȭ1s6@:�	7" �PX�H��R@����׵dUr��[�v�J���4�Z'�)��lĥWL
9��)U����k�u�{��0E�Pg�\�8&4�FUc�t�t��#��-E�B�G��L� ���nh�'N�Q	9����%|����a�m92���Y�h[K&��/$H&�O{4[�!�k{7F[�\�/I�+_��.�~��!���Z��Ѹw�11ū���Y�B��@)�`��hY�h���V��p�� ��1D�����߂�*�ԗOӪ����e��i9`��`:xXP����Ì_�rĎ��׫
�]#
��ʨ9Dj��?Wɋ�ET,L4��wiZ��F<��Ή��v/�Ii;��
��3��f`�7i�r������l �g�`�,Ra�e�ժ���e���ɲ���\y��jj���~:F����]���|m�Tm^��q6���U[1w<�#x�(!����^n;4�d>"�a{���$��%�%p�^��f��ߔI�w�{E�C��k�P-���qf��1޿�Z_�)�7���V���������㶯	�}:?5R�p�o_�W����
�ϼ���%{I�-g�u���,3���;-�qV��ywʲ�gZ#m>w�?�h�^�����'�M:��JU=o��]��:�m.�d<}Y)ҍ|��!���pPn�Ր��;!�*x�(��qzHZ�2|�H����^�mx��]��h~�����>'��)zk���\]�'�@D���e��Љ@K'��Қz��������d�i��d[�N��zn��)Y3���~�9v:���:�?-x��D���h�j`B�򚂘D�^|�ka8G(
�W7:��(,4���>}fw�ˢ�����VQ�!O��k�[�Լ��{�¡xм (� ���ǻN�T�
4��o� bccT�T�Y������s����y0�ЇKp�����)���åO�;��u(���{� �ǆ�n���)��N- �\W���zg@ܵ��ƩJn��+3���kK2�=�;���v˝���I2 �9�`�;P)|J���t���2���R8^��F�	 ~k@'���>��<�ɏ�� Գ�NE��JU�����ӱo�k��ˮ=1%*�[��߀��v9KG�1q�*�Y�.%6LBZ�՟6���O%P���v.�"u�\�[}y�`p�Gk�� ��("�i�x8ą�Y��.�8�7���ea�=0�������%�~[I8��5zm��b�R(�l{ �R���n�W�2�M�e?�-ߢb�B~��m��b@�fѡ�#Z
QSr���b��qb�|0?L�ߢp�$;7a��ɑ��e��aU6��,�Y����8��91`s��E�'h�1�#H��-�q��e=� �"kV��X���A�߳چ�"��faI���;�O!����4z� ��3ksfv-���@�47^��1���ke\R5���e!�vK.#D"w{O�(�Q��b�e���I�O��V(I}ɘϘ|n%���9�b߂�FfF�ʋ��z�{BI��c��!�cw	�?K�r.���Hzl�m��{�C{��6\��6%x@~򀄳�w��UF}��u^֫��S��1;{ˇO���r�a -���9�}Hb%�����:9�&1���?X��7���$�4u����
RHJ�k�r�㧟�#c���aQ��,�]]�4�o]3;^)�<��Wj�X�y��'��<ܥ;+3�D�lc��pDl��B�~Ts�r����6�x���i��9	�)]_*�T*v	1�,o��g�i�3�/��ˏْJn녬�,/+���@�kݭ��$\���-�~<�?��%-5Ɍ8ί
6��V4c������@D�k둚�e�!>�e�M�0�C]�������^B��=5�P�R��FV��,_wI��4�z|����|�����מ�%�0�w���{sD� gi�#�l ����:t���ݑ)�C�<�QTo`ՙ��E���
8l�@<��;4�bXe�����-S7t}Eb�4��3�}Lxo�nZYk��*G�Vo{�%[#��P��/�t����0� `�Z�]�e����:v/t:6�q���H}��AR�8�.NȘMw����z��I�.&��^V�~��u�nr����*�Rh�$^�F�Y;�#�{�8�)?;�}��	M����{����zD����ر��1h��U���R�s�U�ܓ���f����PF�Ӈ�}�@�q���݋��������o�c���Y�"K���`
�j��&q�EVa������{�d���i��5a�� ��
���ͳݓq�:����F7���=E��8�r���4ت+��WF��<�L���i�2��}dt���@m	b?Y{K&3gt�7ؔSq�T�� �K�Я���B���F�'���������/5l����0�ܽ�Xjh���P�<�ƪ�|ST��}��9�;q��=�d]�7�6�Ll����m�� 4ϓ��QL�A�/��Y9dQ�9�5�/-���O��T9�Rhe+>��u����Z%ސ��1+^���ّ�Z�<�&���������P!h�HSDf���}bv�0?�w�A��aWI��5�囀�-
�$�9o+��k>�r�OR���1恓 5�	M���B�����X�v*�nȢz\m-���{*��@��s`4�/a���9M��\����=�� }�Ir�8?_��(�'�n_g��D8p���J���#ϴ�X�~=�D�����=Mf��lp|嵢���Xo�I�\^1�'�U���r�<�#��^�Z�^$+5��V��[�8�òU�I!�Q,gh0G*��⁇�e�3�9!� �p�;p8FJ{G��#/:�S+�6�����d��)�Lo��y��+�-#0��ؼ� ���V�;��K�y˴�8�
��=�PQ�d2r��+���wP4��u%e���]�zt�AF����L�Y�qjFGh���v�?tWn�X\J {���>����Χ[L�ݧ��JD�qp���atp�����xN���9�^�";-�l-��=	|�0�ڄ���㧂�ĵ�ÈN�u���9ԙ}}��H�D�e1����O��A�m���/Ȋz�[�ٚ����$,%շ��G��c���a��B{��D+��pܸ/2��a5QPX�{��v���j��J�B����N.���%x�;��ꉪ�|��}h��!��U�,��x���.OW5� ꢀ��e��s<���{�7ׄW��l��l�XlxVHYEB    fa00    10c0	%(J�-c���}:�G���M|f���&*F�s�X�<��@�^^+�3��������8b�p�$X���g8ĭ��,�iA�FA�ǯ�W�p[1g���`�>�?�W��5�d�� ����G��{�U�˷B�J*qr���Z���dZ���
2ʉil/��9+�����L�H~����HȦ�[��7�w!���<���_����v43�
kڙ|��x��ӼP1$%�J��+"3���݌u�˾.x���WI�3���!��t�9V�Cߞ��sU��b�����fI��,&�%����5������QN��@~���ͳx�Β�Y��Z�Fa�>\���5�Nf�Ʊ�jv)��p�MkV�>�#���;��RC?�t��^���cZ2J`-�� ��7]VM �8U���"��2�?��Ξ�}Ǚ%��s�B5�@;�.dػrS���s<ܽ+7��b̽��#o�|Z.�ɱ�/,�I�E��ed���~�ne[�p��$�v��O�b�M/��R�AO��9|��(ǄK��]��}ϊْ����S@㈎�:���M2�.?�b�����GV�Nױ{�N�#ڛ��c6s�:l"OAtm����}�lN2�A�����ArG��v���:aP��H�R,��~�'m�z�;m����v�1��'�p�A�YA�YVq�gvj�L��]�rf��!\�O�0�x��(�G�)�x�����{x���R��&�o�lA���6�AM(�*��H
P������=�@��a�W
�=�+�&�w�\�rxIU�2:�o0�'�1�/O9h*��T�A��qk*]]�^�;��2�U;x�LX�<�U�
���G�j���4=�������j�v����h/��
���������ma,r�}Hm���M�J~o���D�e�OH@WWK�?t�X��v�aA��ްF]K��z���i��a�t��X���4�gQ�c--�v����ޗ���~KD4��[�9�B�`� k*�h^��c�ar6��?��m��y�0BK�� �礟��%	���X����^gY6��72u�R����0F�Q�d�47��G��ԢRb��>PDe'G��νzWPM�<yD��%P�\|�mX�hH�����J�P��P�$��yL�pK7eV�7JH�e'Eo�&I4ق��oM��l��Z�(~�4_��15�׵�k������uUT4��
Նr:��k����NPD�����؉j+m���1�y�����25�rl3�hI���p�9*<��X�t�s}�¥��~0�~V����4̚�]|T�=�7\jR>����%3�� b�Ͽh�CG�:���ϙ�]�S>��#���DBP�m�tl��6q��:\l/�2��Ύ-�.���3>���9���׽��ey.<`��ģ�<]�B/�D�+iN��'�I�a*:��!��2�┹	W��?���^��Yu�20I/��a��""i�7��U'���]ڱ���(�T��a�H}hR��~{��]���@-�����C���zۮ��3-8��d9rt�zL_f
��}-�W���rL>	a���t�r�����P	3Z�4�@]A�X�I6-�Kq@��v0��^y]'I Tx���^�X!W�`QB77s����Wȫ4��q�9w,Z炐���W�+q{�t� B�[n�� ��ت}��"G�&��Z<�� ����T��C�@ެ�ۿ��}�cðL}��ll�d�U>������PBn!��DI�!H&绖n)�R���_�� E��;��ldb������:�2�O��e:�3�&� e����.�ⶾ|�Q��)@p0���K�F�7/��s�s�B�+�N� Na�wʈ��[�;�)�4uѶz��z�b4ʜ
usmi�[��J�l61��l��|�84��]4SL{�����52Ա�e+�G��RH���w=��v[N(�Z-�R��/�w�J�gG��;�g>^�.�) �}ݽ�ڙK�鍶�k���T�m=�1��+g[Uy|g
#yV��ⳝMM��s����H�v���å,�n� ^K1����R�e�F�AU�z��'�{��JD��{#��k$�.l��,؉�7�|�=��W�����X��&JQX��+��*,�b�%Ȱ���%�1,�#x�>E�|���P���f�r���W/7���L����%m?��!�T�ӭ����=�w����ץC����nfH0�G���� ��|T�~Mo��D7��������$#�}Ͼ�����{ܳU��[G�r���O��*�����(�_��_���!�K�]�x���~W^V�Zv�DZq�X,
U a��-2�f�o0�����u��ʰ(u�\|3���P���o.<�R� p� 7h>�<����A��ک�F��~��>6q�mۆ�~X���V��(ܜ|�+�y�.�*wؖ]�+����v�����{�N��6��l	Ͽ�q��@�6`�!WT5��H��]�x4�P�,k��x��4-�S�������^��������@��q��F�!���(tK�Ok��ǰS�S�D"����sXaT!s���-�@�������(i2̃5'�������>�T�Xdf^��p��ebD'gS��k���� ��~�ڂ3�Eݽ�VԸ�$\���=R�
��1��6�	��>�We��1ˬ�{�s,P�뻔�В,��1.�pM���Ps�m=�U��bL�~��.ڠQ���.9y�35@��	�!
I���E��pl�)\tѹ��j�C�%�)T���1�k��X�tϟ�ԩ�|�NX �[L���uV��+t�cd�'Ff͖n?�4I]%s����M�eK�i֦l+ֵ��2���k�i܄��O9}A�ueX. ��O�� N�/�|�'��.kH���Mk���$.m�~׏"�Լ1#$�uk��I��^w��YN!h[�~?�{��W�X`���'p�͐Kr���0�;�	]�&cp$Z�k�(0���G����pUIl�>� 8e���[�~�^�m�X;#\��n����m���V$���3E4�z��]�Nr��Փ �}���!텒�� ���������
 z#����L�UP9��N�������ysE-ќ"�$E����݂~�[�D�=Xnf���ٵg5��-�e�敼/��쒎Nt�����Tl��Z5Е+UI�VM��������ى�����:�ݠ�ȗM#�u�/.Pߩe �a�	Uz��ݖX� p�.u�^{M���O+فQl��S�"�m���b)�w��G@�	��L(o%�O��8� �2&.d%F�EgM�v�U��m'�~(�EO{����=�.��,QU�$�
��ZaV��_���ƚ�k?�����.�D$����S]�w-;Y�{'�}F�����?�K=`5�(}�ÅC��R��m6,ˌ� ���+�^/_46� ��f&_�|1cX|�y3�&�6��D���������<�����.��f��G�@�@~�4�gt�i"�K�Pz{esV�Nm�Ywp��
�Ck��caz3y�7��.��";�f�&s���徦(�M���8�F�~��u��2���E��vԻ��n�q��#QP`?��vA�f-` d>��Xv섣�F�!�+86�Ə�&����^'��Kr�#>V[��y tx�yHـ�(v5��wF��9T��,����+��K�Gk�]��d���Q��<I���$ⶵ%���~��$C�e������t7cǼ�
X���J������?�d�8Z�r��dD����t4)3!��p�(��zb9�����z;@�\Z�����2����I�3.�e-!�����.E�s$z�#';��s�OJ$�	� SU�a�����I��ՙ�ϼ
��i�S��)��B )��r#3b�w�]Y�6l���<��¢u���>�ɕ�_[@��D��J�TO�P9��²���P��R�wXELVc�ꋟ�z�'���k�C���M
Q��/�
�?@ۂ�cW�����RY
o���	��`�"Y�UyBqͳ���Xd�q�|Z��f�_�0�03|M�UմL&��9iBgʮ�C��� ���$7ϥ�9jU켳g=Nc]/2>֛����+EH��bGZ9HA �%-��*����qIA�"���0�m������%R0��0];����HU�%�v�ف��XlxVHYEB    fa00    1140Q:�r��:%���׼j6�Y='�+h��l�s�����_c|�f.L��D�o���J�_�)�d��@�������x4)RdX�n�%��r��r��J>���E{�t='��zSt�'�gy���@���:�z� �s���LE�bg]	�]2dB�'
�����8N���y��(��n����V�C�b���h�p�A���co�7JR����f6�O���?	���[;����C�1�iylYgUa�y�0���z��ن��|�EM�t��!�Ym�ҽ�Y5P�[��p��KV	f�xJ�#�NAI���bH����iܣ�U� ��0n�Β\���O�/�aQ�q��9J�5d7�0�rV!�%5��Y��{�q��r�/Ї�#���2��r�.��1�Bn��|Wl�Q���<%�q(Zv�����;�����ΓӀ,�w���莢?Y��$� ����JAO�T�:HJ�H:h�j~�ʺ��g�w�YB�D��4����}Zs�7D^
�Bq�&<�+���L�����&B���0%��i�}�nA.{����5Ջ�o[�
*�(��]ĭvF8�����"_�W�v��G��!�$[�/H�;��w�����l�`��&��޼T%.sY���,��\��ǥN61�h��w�9�X��w��w5ӼJ�wQ�\��k(�||��^k=��j��ؔ��la��َ�o�1d*CR��@{O��Bn����oЏJ�_������@��&g���嬺.έRZڡ:���߅�X����DOE.�-�J�Qk�&k��p�z����r�h�����R����i���;مl�(#�9�c���;�gvm�V7�������)>DY���%��K��zp�T�h�
rgepQ϶b8����v.�Ɗ��9C��I��.�e�=T4c�)�n�����=�����E�U�Ǡs�Е[�� x�s�_�몎�w2����m�u��.M�W&����ّ7/A���G��l"�\�2;NҔם�/�k[�gi"�ۑ���� �����]߱D|�h܎��L����%��]�u[ ��?{Oo�߱<�ҫ�F2�j�\�݃�$�����>˄G-�)�KR���'P����8[��F��}��a>d�����_�L���k�R�҅Wf����/zk��,���WTC;�3��D����F�pbv.X��ĺ�TUV�8�s�z��j�O1ST��*�-'7�4�����_Z\Y|��o�Kr.V�*akDg�t�3�"'�o����D�w���R
�}�6q�ؔ�0���F&Ws�)�=��9�}jg�B���)���7V��g#�Gj��.�ԉy�K�a�q�&�e�cn��Pu*gY��ͨ���6˨m���A�������30��1+ox����C�P����6�T��D��S̢���K�v6�����˙�nb��J�<ۖ�:��³����oxj�^��N8�Ñ�cbf��gWK�".B����Cҏ׊��[ѭ�wz5eR��)FA���IH*\��a�B������o�vZ�ۺ"�y�{22S[c��G��n��H�Su1��5�!����� ��@��h#n��L�Y��4�g�5��q+���G�xV?��QOeֺYH�v��j�9ƳA���#��E+�����Tl/�#`��K(� \w�T�KUj(���	����;Qe��N�Lu�w-�����߂
�05�X�`�"��k%�.�c�����,��1���،ށ�mi���?���6����Ž8~�/��Ll]t����v�«V���ne��Q��_P9��RRA���n�wokC̭>�z��I��HĦ�|�?� Av���cF���JJy����7��?��q�����)7�Ľ����*��|���bZ�wD5U!
A�'�O�0j`Y�T3D���3кz6���gߏ�Bw���,��߮6��#��z��5&k��O�|Lt�z<ͼnS��Sx;2w�R^��G�U�]�ߕ�I�Y�?����+��u��P��4�4�{�57CԌ�ܜ��P ��7���s�|�3�ڨ��R������<��ȭ.��yf��`vx[�^N7�8G����q�#�
֞������cV�;�t]��1�ݹ�5��-Sщw�VZ��!#�f���c��&�� �%ۧu�@�O�Q�ߵ�c��A�m��=�g&��F��/�V(Y��/ɣ=��㢹
=�1���3xq�+*���Z�9���5{�u#�0��z����&�i��k�k5���Q�򥃉�/�]ē8�)Y�Jh���N��1@�v�Ѡ��-K 9v��zTo����mw�8��ww�X M����xh�ơ�∭���&ۮ��M�Ook�`� M���L�03
�ʊ���8���E��i�Sd���N��;LeqLF(�"��Y����$N٤���Ϧ�	�"�ɔ�T���W�6���&򷁙��x{����e�w<��q�(���񆰣�J� �uҴ�u0}w*O��!�Q?��Ô��RFN��u��IY���\��Ñ��h�F�">���u)$�e��QFH�7�`1���N�8'U��7�:�2�q�!��q6�[m�������)�?�B�Q��4�v�gt���-j\x>��S�H���e~6)fx��G��%��-�H����-������e��#�ʈ{�����w�y8}����-��K-�Ha�81{�u�4�N�i�gƟc��gH��ID4��ͩ@��ɖ٧��r
����7 o��U� ��5-?�_5�#��l�:(6��U98��^��B�<�5@LKvf��*%�x�V��Q;uA4<� �>��P�F����yl�I����M0ߎ�\~�K�x H{;G�r/%bO�ye���s�,��Vf��w��=�r�-gݲ���?���<]��.:�������K�����Qp	T�@�Oy������33�Q��C����%Q2���Oh{��%��R�R$x��)�wm�qj��'À򺈮��K99�Ck��6}!����:`����!rIC?�K����@�feNI��u��딉�;Y����ld���'��u&`��Mn����o�na��������$M{�L��u���M	�sVoq7n��TnJ�Z��쳴�-f\^_�*���#��L}E�S�u�@ه�
���`4T�W�j%J��Na4g�u�e6�{�,��tF�� V�?@&�g�=QU���rd���_�(8�a�'�RU�|eM3F����;��֒m�� y�@K�j�h�0�{.z��{d�]*0^��G���#��r��~9a�h���$ȧ�[��DI>���n�a��g�c|�7�r#��o��6�Q$o���8�O�$&s��h����;	�q��.��`h�:�8�#T>ϐ�ť�u!a����<�V4��]C��iN���2ӔpS�O�E8�3�Zo������@���Ue��w�e�ʀ6����i>�nQ�dPR�qRp�Q
������퇾��iv���ث���;]c��H^l-�W�E�J� ��5�O[hG�b`4-1S8�_���n����K��l��t���n��"�;[�>��2��\����wl>���V��H�Њ�ƔM<��D�F����<!�qQ�fR4�S3�ۏM�P��5~�BrC#��#j2�v_�qZ$S)"s�����`�rU˞��/R������2y�|w��,�G���!.�Gp���RL���\�&snV��"~�A�+w�u
���F��.y,jJ�nE�"����Vs�������/�Č{7����"���O�h����u�_0'tw�����Ǘ�z_���z��Kkq��=ֻ����W�$�*���As#\��������Z9> rM�|L�05 �����=����Z�h U�>���Oh>-���?����Zo�ߘy����T��o��,�-�Y�r@��꙲�H[�T$���썧���ҹ�*@����h�Rx;V�!��c���3/g	���>�\��l���D,�Cj��}{�u:���HD$���8��<�	4E�om�#Y`p�k�O�Y`����+,��@C1���Nd��dms���L�>BSS�h��G��9�Лr%�c�`�T��o���̨��-Y�#c2aj#���a�I�-6]�c�	������V���̂9��H���y�`C��.�"���^�"ft��'�t�l�J���F��U�1��
��"�%=�y��<>�]���|� H(3����-�_U-ت�{'��.��"{%�c
��#�'��I�5�|&�o8T�]��{�Z0P�����Ġ��ф�Kv�ߪZ�(
k���e� �``�>8XlxVHYEB    fa00    12e0j+��7-u2��Q��';�b`IM|�'�J2nq̓�	ß|~ҟ�z���MF��h��a���C�����f4pt ľpK��z�}�{ё�b �V�h�nH2b֫!,9-9"cΛW
B�� �ǡ�T�8\0�1���-`��J/��R뮪�x%���2�!"�I��C��<V.�V�q�~i�����/�pǂ0�e
3�����>���֝�x��R��7�uz<�T�dkj�7��M��|M�(��6��텥��Z���G�@�X���uV�u��
�����k�<A=��#����0� �.b��$p�>�Hw�n�����dՃ���W&䫱^!徦�p�Q�;��ߎ[[�cceO	̂l�T�Izk�$��O���!�0�W-�4� �'^��%Ylx\\O��3�;5�y㫙Y��k�kǲV�Y4`ǿ�>�;z�3���#�#�uh�h��?.�	�9�>���=�E��*|]��Ko���� ��$�޾O�pm�TPR��Ƶr�;v���1�np�Qu� ���S(��,p�lC}��LJ��'/�0*��5����תT�? ����ߠ$���y�i�@4���^y#D����rC���|w{�ͮ��L���і!ܒR́�i:U�ZB�6�h�x��iCj��}�&Z� Hj!2�h���_X��r����~7���U"N$�fI!��ZC X8C��ho��U�5�n���B^]�����ʒ�i:2��a'A����QV��I&�<��������lK�9p$��r8�_,8svd�{�q���!�rZ>�,�a18K�岅�`����ђw��:�dm�� �Q��[S��a	A0=T�ʌ�)p������ʨq)��Q9i77��*��%Jh��Iì���Ŕ�Z�Jx ���2Qzۧtf�yّ��SI,}�E
Jv[k�M-����ap����3��p������@ 2�����,�}*i�j��&�m��R���{R�"����T� e�9',�})��ȇM��99P�Ey{ڒ����e�7\n�,��Q��D�S��9�%��k^JD\�������T��+б�Ys~Ɓ�[Đ)|.�һ����po����ھv#y����>-#Ƙʽ��U�-�!�u}�w<�����������,l�f�8�q,fq�ٔ����K�>�
4������(H�6rT9KG����-@u+� �	JVy!�t8%�?�|SH��-l>gH9i�0��I�������x��y[�89�q$M�,,ɤj���R�7n3Cҷ���~�e��ǫ�t�l3���.����%k��Z*`��HO�75�ԉ�����	�q�' �\�����ٶ�
�fd�Eo��Zz_-�9��KC_�ܗfZ�;y+���̦���|7�=|�����;�6���&.�'g��s(��i��6��-���I���۔�^�egKr�'�\�����[LC��Z����nS���0�S�I���D7w��lm�}J���w��A���]}�� �M[m�C)��"��AΤ�䯅H�p^ɾ�^�-�`�Aܔ��	����x�겮ë	��q�嘶h-O�Q��U�/ty��<�,��e� ���e��Nk~Io
����il�Q9`��/���i_��pz:��lek��y�7M�����'�J�av?4�v�Tfa���X`.�]I�X�j_��4����w]��*���k�m��/���W�`�,�E��#�aʡ���l=��n݈*��~/�-з-�K���G�Q������SaeK
Wec"-�VlES��X���9�tu�Ndy���YE��?Z��?��P�H5�j���a.�$g��0]��\I�G�'K���Z6W5^Ti�]n��8L�f�īB�۸	��JL�h֢�E0T
�
�&�}����3�>�+|F`���M�8޷��0a����\��j��V�S�rd��P�E��o8~ �j���!J���7�Hj�r�1�"a5��͋|�R�����B�/њ��{Y�ŵn�"��K�dZ��:�?��KM.K�nrb�]{ ��אdȄ�"b������&��4ɒ�i�B$��c����9;���9d�s �!?@~I)��R�LR�P��9��貎ſ,q��S�����y�eĝ��E��w�rض.��O�u�`e�)U�j:�q�e궣y�5��ꠋ�v*��f��K۽3`ޕ�^��I�b��l��ߌ����'�/�D�in��T�SUN�z� A�e��q�8�����U(��||�m�7��8��V��ŋ�:�V�q�^����j!��&�||�*͢0ã/���K�������"�MJ�#�`�7�q�֪��&'a�]sk�ӧg~F?�@P�.�S��8|�3�1��Y�Z���6D7�_m��e�`vı��j�~���,��;�����C�j�]W�o$�!�;~aY.��݌�N+1]H!�=��"X)�c�;*F���=lc���Oܠ���{�WJ�Mʉ�����i0��c������l�f8�ӆ{���l�>؄�%��ns�)ks����:�U�yBχn����-�Wl�	2��0<�v�%Ș��N\7�G+HZU�Cw8,��z<�8����}�/�m~3����mVD/�ػ*�b�Љ�E�@},?7G�W�v���?�]1X]�1�i\
[[�i�h�
��D�D��/v��9{��ӷ�Sx�����{���\����)�ge4�v��~.�0�H3R،�4�����v��ǈ�})��ü����oӔ����H+����f����:�3,��}���;@!��?d߼_[w�*���~$X���j�πsŔ5��W�X[���n�J)��Z�lA]_F�D�i��,6�_��Ȋ�j����o� �-p�����?!4��R�,Ȕ���oɩ�X �d�j/�SA�&�-b����š-�r�U�j����˹���И`׍�W����G�̗��:^����a6��O�Q�Z�[���s�3:|4����<ip� 2g�>���_��4��3�S����i�SF��|�uw�YM�N�&��ɿ+�:=w�Kv��]n\�E�#7��[O��.�?�����[��D~�Q�������ʇ�>ߵL���[�ٹ���Z��������k�o˴/����AP]�Ϸi��[@�_#�2biFQ��p+:(���4����e��=���"��L@i���CH��CN�jƍ���#��<T֧v�E�yҹG�1�^["������O�,5R�DY���[�}�U���yŰ�$ ��7y���5�Y�����&��g4l��;�&�j&���|��,NfW�"�_��&�ܖZo�\ͱ��H��w��A4⳩O�7�A�
����[�I �sM�_�O�=�o���L��R��+�y-8�N�+\�U'�	�:�v���ؐ��m��U�-��o���Ǝ.H�))$[	��_�g	A�0#d
,F/#Dv�L*�7�H;���)���A	j#�h�!𿧒�iq�|G�d��~e�=���%�'A���{ז{_���|�ʀ�CK��>WQu�x4�HY�����^
������uD.wL�I���9q)�r�Y�U���$���դ�\ٮތ���3Ul�ߛ�LG`澣1�q�m�ڭ��W�R*Ȇ]7@ȷ.A�x[jVQ_[Ƀ�6�,�n��@p7��pz��Җ�Y͌�>>��dMJ1��&_��.���!�~x��*Lw�?�����>l���ʸ�ƌ�P��{Xt��ȫj��+o8X�l�(�"3n��MQ���|9��	?(|X;`��\���
��e<I�td�0px��]��x|fU�pN�q7�v;���w|������-�AF�V�KPeL�j�%�j8P��f�]N}Wip�B~�P��X7[L �?,٬r��yn�V8N *�K]o��J00�o)�gr:��%�;�2��������#��cU�O;��(��zthD��{e��~��a��~��A.Q�rЅL�h0�sW<�����R����w�(�t�z��mЕ�6r,<D��*�p�1K� ;�u'8Bս%n@l����,��k�i�ҰB�ҝ�.���x\ҟ6i ������K��n%��D[����?���Z��/��@��'�`����6k�1������@��M.��[*��0�Ñc�&�Y`1��Q+&�����p�5�6��jM��H9}����2W}�}�ӏ0��Q�Ͼ�H�,�lf���#��e��(�u54�6��
6 ���D�X�x覸�N|��P��v�.���C�>�-�Ă�E�܉=��H��̳o�K��Z��������D̮��[�b�����xA*�����u~�'g��=rP��e��!G��7�����j�f\��X.Z���=��K_q	���6.��z��|�*N��}7��\��w���b|���G��J��Ji����q���?*��t�`(z�VI;�}�r����lz��`C�k��;\>�?�BIG�!�?{��9@��[j$B!�)=�5緉���<�Ӯ�=j�1��ƅp���'�:P)F�]�5��
>�q���|�s�H�_�~�,�f��~�#��9������])=�U�4
��tg�TB����5�Xs�}4�>��BW��$�c�B�#�@�ˁ8����{�C�)��	�+�j�p��q�Z?�&3�{(�˹T��ki6�"�J�x[Ң/��ts���W��:w�鶆	��5XlxVHYEB    fa00     f50�48��y�A4ɹܭiǡ=oewB���h�b	`K���j�.���J%�t2#��0;���[/�����l��2l�hZD9��b���׾6U�ie�	4�R`�VE���f��uE4X�3��Fs-��ص�3�o�!o#D�(���^��/��YG���mtw���^r�.c�v_��H(%��Ȅ1�>�ߵxLO��uLu��y�;U�W��:a�A��O��j�����;'��.�R��5~/UekI)ﳝ>�e����[=�|���u���wU|})��zoդ����?����u������ ̎�W5�םE���i&���D��c�qo��� �րs7X�;��G��ol#�^v?�5\$�`b3?
7�$5A���_џ)^QYjK����S #���"/9�4_�t^H�}=�L����L��svʓ�pևs0�w��U:�2ӎq��g䵎�+��/��u�����`�/�@������$y�� �|z�n�;Ņ*Ŕ��W�q�ޱ��.���<3K��ץ�������y��-�5U�� �0� �w��Od���9b5j5	�
�v��}����̢k:�+�����*�-L�z��U�J�T�ǀOU�Т���t���`�2ASp�G���/$�#��,�c�㙁���F��B;�C.f?N�'ج�`8�7��=M��ݏ��Ƶql��Q�Хn��I���/�Fvq��Y7 aȉ[DV��i�+ly[ ֿ��OXK zpp�'hՅo<}>4b-Lc��!�s}"58Cb�C�z���qHݜ�=R�#����4�/�sk�rYB#�$˳�N* ����aYy�&��� �̽
Վc� 6���%&��_k0e��?C��n�+���#��_�?�VcGw8�JR��}伙Ϡ�9�P.��s߷A�3������}t�KtZ��	����k]|Ny�_�p�N�P"�̱�xw4��y�5�)?ͮ���@Г;�&���d�(���;\��m�M�70��^Y���D��B �;4����{{�U�A�������R��?���C��E�Ŀ�>|r�(��QR�Ǣ2ct��������n�i��a��	��k�w]�����˫�`Ы�erw�@ͨ�s�rՊ�w���Ś�h2���7��ݽ{���."�l���X��E1�϶��� v��H�m��0�<��f�G`2�� �atV�b1&"�v��p� c�.���O�˒�i� !�zwK�ѱ'Y��*�	�MV����e��i���d����rDs^� �|��w\}��r�aca��勤V�ʥ�2{�:9���=R@۴�C��"&F��K�YǾ�B�+��b�"���x�L�Ŗ5��%*��JH�c=%{�Û!S����y�ux1�������i������pK����ש�#��dT�ڼ<�Ԧ��ٗV�J����e���� ����_�{xI�n���'���������V��<04�-�x��~�������0*ʍE��\1�i1#@�C�6yv��\���ͅ��d��D�m�z�;�CFM���L�#��CK��W|����N\�^��[>��7l����]'���O���Jju���5#�87�,�V��L��S9�E�4{#�]
b�g����H��F�������Zw������FO��/�q��DV���&�R3uٞG=��@��E�8�Ľí�%�����pe��0��N���æw�RӁBB�a���o8@�\s?��U�@b�<N�SH����_S��D7���1�R'#�x�ߏ���>�rK�5#�'d�[�S���v�"�r
��i������:~�a���>;Y6������� Cz%�"��e%��W���z	��(+��MO�?.	`��|�/h49ڔ�ݩ���C����\Q�Kqݢx�s��#颁�/����}�=�.�/01ظ�B�컾�c����0*���9� �7��ȳ�|�
������e�RO���tƇ�F�l��6W��{,,��o��U����_c	`�F/7��~�������d�F���.2�}��UP:���[����=�����R��1����}|�����#f���H8Y���ë� �I�8W�x}$9$$�G�<�y)@_qm��=�~��v�F���0�Ɨ��>���=I�Կ�5���u�݋�P<������PT�j���릳_G��ݲ�_�$��b3<����N����q+i�S(l/�?h�ڎ�.��8Y�ҙD0V�2�A\&�2�����K��P��'lu��#9���:��ˤm78�[E�r�ȁ Z���ú3���
w�O�{�Fs�Uo>d��Fp�B����vH�o�_��<)����$�$��4_Ĭ��͗~/=+��X�b�u��Qéc&&�a��)^�e%՞].�p1'pN�j�`�R���:~����E&�2�̫���̎�v��M��YgT��R���������k��9���#������4{��^�r}M�d�� �����7�:I6-�N�3��,j6C�3�""G|�[¿�A� @?W�a�$ W/69Y(�2G�Et^��>��ܲn���vH�-���~5�M%�JPH֬��b_���sKh5㯭�G3��%d^�`�g���ɷ��sqA���[�pV	�*n���O��+Wbw�S���<"��r�t�ﶊ�Ԧ?	�9Ae�6���@X��*U�.I)�,8;��G'���Vc}ݾʕnձ�-x���9����ЗTx<�VG�K�%��T��3Mqjh#}xm��3�!�Xr� �_���U<�;�X�)�����j�t6�LB��7����m��􊟞��ɲ�6φZ�ŏ�6�y�_��,T\Ǝ���� m��ƌ�[�#�y��Kli>/N��ߊ	ż@p\C�,E��J��X���G�Ӷ�'�۝�C���ҿ��v��4Ic��чuV�I���O��+����oA���X�r��ھ�����Y��bƭ�>h`��\�9���z��7�^�o�[�G״�l�h�0��!�Z�hp�Q�Y�lShpIթ���_3H�4�Y�t�lH�`�;��C�m,���v��r��F���a���.����J��m��Wuo~�΁:�#��K��+�8����,�]V�s_�vH���ISZ�xTʍbH�G��\�7��c�)��-[~vN!�YW�,���jx��c�_'�<��@�S"�|	�S�/�nʦ��ȩ�C�̇�r�߱�r1�48N�E��!�����T�;^�i7����I"y����Y�1�H�0�6����Te)Q��^�=԰Ѻ����e��`5��\�- "ԍI�,���M�Q}k����/�k��p�˦���M��%�h����izS7'�h&x����0?��4�L��W���%��ܨ�u%`�Qxx�.P��u��|[��7��
�w��f��P=J�}|�`6��5y4ےl��r�j2xf��"&q�@�N]��������m�;�t���q������[c-��ÖX1ѳ�����G}��E�]�[w@���6������o��@����I�&M�:'�F�eD2��xfė�|=u���+�pvLX܏�-��F������!�:C��֒E��v����߂x�-@���h�@��CHV�+�:��:��q�*��V���D�A��ܩ�a�V�"�z�������x?�
T��P���� y>n�[=c�O�_�ߵc��kՆ�s�OG�C^cg��lZK+s_�1�{�m�uW`u0��]'�ɼqiDM�"�d-���Cn�&!��idzR�9�6���M�0w�X�v��-Iuɨ��r��s�P+/G.���Pe�rXlxVHYEB    7273     560��w.A�c�-�.GT�Q��C#��mOC =�Rbd�H3���@?V�ꚦ����RO�5�}N�N��p#u��^�q�A�z6	y���!�]n1I�|a�t��, �	K����й����㳓�T�y4K̄���G��ÿ6N�S�+���`�W�	Y��* �G(o��w50\[>b9��v������7LH�@kq��Q���	��P!8^c�z�nxX؇�iM���/ �M�𦶎�x�D흛�:ة̉�r�4��xdw��L1(ٻ4da��|�Y�t6E��2���������CA�'�~2p|e.�-��iw�n#nw�c�+_�<�'(}���ּ�V���c������O6r��j���\�I����Xl8nE�h;�Ӎ�65��xj���ª�ZE�3Ee���@���NY��m���aD��ZWZ�e��/i�#�C%��Q�rO�{rB���b4˶�N�h�T!��z�W.^�c*/v ��y�З�\N���[�ܹ��XR8d��EF����O�o9؃S�Xh�ō}��pW��E=�%r���L�_%k���L�Fs�e^e���n7Fg찀+-lߗ�eH��[5��Y*ܖ^(��|��
�c=���#	�s�0�,�Í�Mjr�`�)iIL�zu^�1��v���C c
&�FF��ؔ�%�$��#N8�!�����?4a�3�Wܣ��MM"EC6��� ;�����y?��P��"6�G��y��FQ�O�ut8���[.�>N�M����P�ā��]�d$��Or^�|v�D@@"���ᜥ��7wd����@6�AW�`����m)�g���u�1�(���&;�a��֥��Xٶޏ�c�Z����ya���}�&�P�jjȳ���'�� ����0J}���!��"�E�Z3�0��kE�=����?�n{����U��s�S��xji�5ɲ��Db*�a��Yh�.%���p�A�:�$b� �V�ؕ�(�H�����'�LO\*n�/�[/2�<7ጐ�Wa�6jUk\ m�]DdNE���N���E�;;rG`�}�]c����N]�k3x�Z���;�٢�	�)���o��A����q�.=���%�\��;���_KjQ�	\�F���K�0I��6��*��(�p8��1��J��ڮrb�<�Zv��8y��� 6L�����EW'97���`k�k������p�b�|J�!��wX�MQ���d��P]-�M�e��.B�1|]��3�K��WJ�W�4C4y�m���`��XC�f�ȷ���o��I<��xS7����Wӫ<YUz!�#�@k���>���� \��Yy�ԁ����~��y���h�-��ot