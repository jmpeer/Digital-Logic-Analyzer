XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/����ݎ��z����#��̐�.J>[�TI���U�]��=����ǉ��/H�&>������n��s�M�&`��W]����a��<��3=��6��6FU���sۊ 
&jg.#@��<O7�.�[i9\{����.$���"��n
ȃw���Ea��$�>��m�ca�~m���T{�Q˟ښIt5����Q"FX���{;� ���*�	�Wn-��DB�0��^$��C�Dr:~��)%�F�ܽ�'���WUK��y��?����s��O�~�;�53H���z5�~�.Y�,��1�Sr��40�������+Z��ė|��
���#�������;-�U}��sL��l��I�{�cWY�����X;��^h�/c4K��!0���ר��e	n�i�81
��I��J,Ko�<��S"��(�5}�!�����cZ	�aF�9~;�8�|��p�A\�ͮ�D1�Ր�8���vk4�)�3���%�(a�gl�]E$�[Re	�>�(�tN�h!�0�!6���OV8�
"��6�vaMN��[�'g��C�ٌ�cޓ)H�K���_��o�Nל5�t����Zj�����k߶�e&4̣-��56Qݺ�����h�I;7�V�_�R�+�OV~�E�ݯ�-�
ԅfK��R�b���:�(V�U[rT�Kr�j&����X�V�rF(�}v�������Qq<�:�1���	��<���1�P�A�QL38��S�"$|��M%�#rDΈ���MGjì�><��[�z�XlxVHYEB    fa00    2260�%z"��L(Hw�ʗ]1%J)#.�M:O񙻐zsl��1Vf;in��8ظG#�ݒoU?�EZ��j�o�xDuW8�G2��tm��s6a��[���k`_�wrn{�V����<{���V� ��m6���	�S?"(9�J���/Lt�v�rM0�%8�g���k�[4�sH.U���t�@��Ns��1$|�	����}z���k�&p-��K��%.�#�w������ײ�B�����w	J�Ee�˨�mл�'_��醎��/������9)������nw���EV�5�[�V�@,�[��x�d��6�����؀���23�c]���R����H�����GD�v��᏿��eV�� ��`M�@.�R*���5M���y5/1�ZL�9!��Ǹ�nY��+�fLy=�.�+�""��7&9��_^5H��nG:��T���=G�b�4���[���v.g�t�e׌��~��J�n��=�����ɺZ-�9��
����,�"���|h�z�?Y��)�y
)J��'��x�}d��IVM:��P~��Dt��>����Z���xju��=���]��u.��*��R(�-��n��ץ,��g��8�x?�eX�i���O� �Tn�H��_"+�L�1�]���\�Z߹ns37�W��Ytt��ّ֟#M�ݬTݿ :���{��F1H��-�]
�_�f�=�{8�}��+�Z�G�H�H#t�c�%i�'�����j����g��
S�9�.;#��~&���X:�+���z�*��!:0���ı���`��scSo84GYI�!^�ݭ�)2v�b��7����h"�\o=��Vи{�l�K�q�_�w@�����Q�l��an��(��r_��ZeK*�l��5o�m �?Eq����Ьr��r}���)'�Bl��G�0�4"�����'�����Ɗ���Q���R����zu<P���[����1���d��\Ү|V����6(�4��b:#�U/¸�j�\�	���;���Z��}����J�e|��g8��k^���_�f�?�I�Ly/��o6$}��N/���Ǝ^���&����-S��h�}c�̴DӠtg�a�!j�6�G"��6�doI: bD���٨�P3�C!���.������ �teUf�.I��[�z��WZ�ǌ�wLG�5���#l��L��<p	�i�J�[to�,Ū��'��#�o�/x
�z>	���,O�c�
~^�����3���X�g�7�x����<�����i�q�_e�ş>�{�?U�j�^������E6N��@<���rnA��x��LZP�}�U�5|q�~���ݻ9H4
ch=�[�XF��B�.�<s^M���xAIt (=8�FtX��j���^r��`ɟ��7D��p�b)7�$��zA�� D�Q���T��w�F�F���q�:�X�o��c�f�{�+=&d�!���=p�5x���Y����	H����a7���JK+�뭾��D�D��T¡�`f�'Jq��65�@�M�_w�/M�G}�J�=��	��)lʳi�pл���ğ�tW~�8Ù��)�V��s�x����u�.+r��k<� ܣb��	��=�����rQ���8S�!Q� 6�.��Pm��w)�j���U(�׀Q�6�>�dWC\�����E��	#5�V8�~p�P��Q����K�n����7I*�B�?��_�,�=��Ck��K����
ѕ�οP��n0Y��`���S�z��ǇE	�����7<|�"=��ɤR�iѩ㒄�WY����ظ�]�| +�5��4�����Q�k�����:�?0�\��Q�d!���y�'���~�S&9/z�j}�eR6���:-�~1}�V��V�������N�_g�0�h� I7P��XRoQ�HU��r.�zM�f@�a���s��X�/��z�w��6�E�����&��WR�ט� �dWN��9�/۸Z�=7�OF[!wt���VC��6�� �8��MK����6s���_�E��i�]0�n?���:pU�t����Sh<�JNK���(ҥBe�ը[�H�����aD-9DsP��A�=_U���>�@���h�NJ]F��$+���ФAg4zF?d���CK� *�=����g�<
�W�H-�P���d,����	<sN\mӫ:�QL'�m�Ez�7sA��0�6���K+D�+G9�O�(�vx�1g��7`�{'l���K��[���-^YW�<O�ם��W"gՉ�>uҤj���x<�"c�=i(�#�q�$*ϊy�.�"���y�y��p����c"��a���A����lUe��hQ=��2����9M��1�YEfދ|��<+�v���+���7UƁM������`���P�l�!	�L�hR>=,�|45.Y$����:���,����Gz�8��'���L��E�,��+�|��G5���[L����l�6�Z��l
1��US���Át\����7�v���)
��$�O
W�<���qX�?+T
F���S�>��k��V����;W�S��[p�c��Ք��O�mY_9��{�]%�R<6׭w6�$��y+�eQHgc�H2��ߩ�)����=I���/�i��b(��=2dk:ͻ\�~C��{��S�X�����U��pRE�p���[���:,�����6���J(|������V~�K�=<oW�y��X�{�^��抺	��Ӫ|-(!�9w�]�������>ju�h}�'ɲ����[¼�Z�P��ޏ��{?2foYy�FĔ6�HQ�r��0Ύ��Q�D�n��m��R75%�qu	$CT-B�6��;mz���7+z�ݷ�ڇ���  0_���OS1��u�,�+R~�nÖ���א����(y��3��3�O=�{ m�ͦ�=��v=�a���1z��g3�I����G�m���B�����1/�*�W�	  F���[��|E Sh�V`�?�o�|[P[ʘ�y~���ST(���xN�78�I����5`Y�p�PW��G*��U��z�a�&��^F�s9��#ڻ��^���L�+��[<5�;�Pj���V7�E�ȿ�ӝ#=�(6�^_����$+���d�m�+�ڨ23�q��
�WA�ѼI���#��;zX��HU���n��гtJ�V
��ݏD��X���x��gVR���$!����[2UcKK��a�y�˪q�/Gv�,$�v̨�;�G	�NV��u[�;��ъ���خ/�,��¢s*5&~!��K����]=���ܶ}{v{,�YG�d/�r=>�r�H`)����J��v3�@Di�A��k��ܘ����u.���ZS
��J.u1��^j��\���?G1�ٮ=}K֖�RS�v2�l/�M$WF+�	��
�]�]��E�_� �b�X��:^3gSb��"�t�������y� ����)]�����]F��&��I��i~+Z�_*�SN���{��K+�6Y��������9���lQ��Mc��t���{��|1�[�L��Vϗ��B�8�ECr�n�g*����]�*�X����BI��,�W�e�۲�=�����Y��2b�w�{�9I7��\�mN���u7�e�ld��[ #��%J�H	-/rِÿ�4ʷ���Dy&o�����:7*�>� AR?��O�'���m1^Q�s�kگLL�ho�*ߔa����K��sɖZ�t6@�i�[%&;�#��Pa�}5�`'���d��Z4:�x6��ZL�@�|�<�2�M�E��ǒt��y~��	q>*?���
a Pũ,i,�&��o����/�_��� �:�`ܫ�sjlE�x%~,��i�]0���F�"��Pą/dBb�-���j�'s�yM)��5��ۉt#���@��Od\���CO=�6|]$���<8lE%�ߊ+-�F��,K6�3��Njx����8M��}�E�#+�� �6��|��H�G������<G����0#q�ڢـL����p��+����&���q/����Nt�;���@u'`"������1`�',��9���.\}��t��<����0���_���W�U��� �q��k�e5�����|��[�2
����@�,&��wj��o���Z#'�
M @;k��F!KI'�Iq"�d�yT�R��KNLt����]��˨�$;�չ��:u d� �c������zi{H'@�� w���CY������0z:$�Jo��<m���݆�����y���n�߰z. fW�r�˾׬��H����{X��"�����$C�ԝ��ܭʦR�,d�(߶Э�I���Ќ{M]��ii}_e�ͥ�7'���yQ����a�)�C7$ZI/]**z��)�A���:n�^P�f�w �:����������`qю$��m�����:�"��Z��+�5nԪ��76P��P�&*�g��Zte)M�Em��0�X�5�W��ه��?AS2�ń'J�����A�j�aFE�G\{�`wYF�"�:U����I��dDe�ŵ�`���D|NY4�B?�B���A���<��$�F\K�A�����0P+w��a4_ϙ�Jo��V����MXkˢ<	�P���Eb��ҟ��̳��#�9���Tq�pS�j8����ʈY�]�I`,���+���ꤚ�A�L���@͞�Jt�Wɛ�I|Q��8I\R&q�����F��k�vE���X��4J�'ڎ��������!;�hIy}W�;�)�+�h�6�w��!�����DD�{�Cr�6����(�-�[zb�8tޑ�P�����#'ޭ�����ص�5�s�8Cےn"�C��k8�xZf�PJ���jD�3����?��~z^iq�����~��C�i�xO'��x?&@�Jj��P��4ω��q ��%�A���"��ͼ�Oa�O�˼�/K��=�<�n��`�?s�뀧��]b�� d_1�5�ᖮQ6���S���P�� ��U�����r-�Bݻ���TN�#,������ހ����g*]���vx��^p��)k�������s*;��3tR�/Ab���k��|_��b͚��9�����En��Ŧ���+��x�x�᪾'�:y^c&E|["Y��0S�d��m]K�#	��
@E'�������[� í����<��;~9����=���T�0�p�U���*j͒��X��ƌ�x�y^�w"��j������ȹ�w��}�HC!�F^���/ofR�Đ��U��& �:C&���I]6��� ��}�@	m�^ǥ���LY":u2�z�	`�T�W�	���{"���,.����|��b?�̱z��zp��F�����D�E5B*�>�#X��mQ�(&��Q��xsy�鴗�X��B��Rk%���v#
>W
��|&�!�����g�2!z����YLP�S0m�lr^ž��RH��o�Z�4y{�xq:" �Z�.��佇aC��-!�bT��I�uT���#E��(K"�9���61(��}�I��<�<�n�H�7վ�.�؜��$� ��B�!V��J@WK�wi��Г�07�w���+)~����b�sc�+j���N���"�`J���ӕ���z8d�z�E�G��w���^,��?�VЋ��a����G,7�����%*���\~��v"�;��]�r�K������ ����:��������xi�fJuV9i���}I����ȳ�k�_J�AG�
V k������s�A�ڝ�s��w�*�+g���{IG���0���[00�@Ciu5�5ا�o������h��}��p��t����b�}���e~Į.�ߴ��h_�N�,�5���F�@��a��#�dZʽpA�F�@
ˀ
�O�Fj���RP'�I<]/�=���,� �N%�v�����rRvc�Yp|�jE�Ͷ~�D�&��U��X,boz2l�U,����}ʚQ���6��sק$���]l�ԭ#�1d���W�u�b]�����C��=.���>Y\s�)ɘ]{Qp0ҫ�l\���i,�ȧ�����2N��S��{��٠S1$���c�������+ΩPS�i�(��$�U��Q���s.����"\�$������b���|�fo�!�9#�ì��*��t<d}�Zh�;���t��ڈ*�A�[�F�� �S�S����
/b�ܝ� �<$L�Y��?˟qU��WFz���(�gA8���d��iJ�#�����	�1����$��!������%O-H>�܉��}�w��a��̮�_V�ۊ����.j}��A�eE%�b���_�
w���_|g�ɣ% �"��孀6Deɋt�=i$�Q�*fF<�f�F��h���5H��묎�l��K6�]~Z`���W��ƫ�{�̏0�0���W'h��t�q� ��D�'S+�2oL�,_�wY:��Ĩ����t�p����Ǉ�*�&�[v����Ӭ	�75��iF�Z�|ۍپv(��I��@Y����ik������\����Ď�NC�Mo%�E0&g�f������Ct#��7t˅�IwI2���9l����B|,���P�5�IZ�(MgܯUmJr \����VW��&�N��e�7�He�gV^��R�S"#33��I�4/B���S�f6�(0A�Hy����J�ᏸ�|������O?%�-��?qV�\�=1�|��BM��}��j�����?^O[A8GA䃇��+��'U/9��7,G7�O�~�����<�D6� Z�@=Q��0FwtD Q@��J�<C��!p���d�W���t1�D.�}*���P�^.�](��b�y�B��*ude�	U��PxEϋ�\��67��s$@^����!�%b8�#z�N��#�ݯd���!)�����6���X�&z$!�F�ԓT���Z���u�H��:����{l\a��W�j?�.��
yemR��R�EO���uѬk�6'y_�21��I���̞�u.$A��u�+��W�_Y���V�cJ/bs�����b��1p����񅏇a�沵`�*m5t��";(���4��fݍ����r���I���r8��WOS��
_�"t/^�D���W���B� v:�B���~�(D�-��L�z l��1�ͻ�U���?aCt�5`[��Jh�V��N�?�F���%����F`��8f�y
ˣ�>c������5�E�o�U�k���ûO4sT�L�u-`e�o�$�׺y)9�Cy{$�y4�N�0+�#	��|xp'�ڂ]u��@kJ�k:�;�ȟ���Y��~��0�N�`��p�r*L�� �wq�v$ ��!L��(k��u�@^�6�GYF'P�d�8,�� �AO�p��偒$�"^W�9;
�u�R���w�y;2p��1͜�![@f�vE��=|o\��yT��į*�X�X@�!Da� H鬎��%u���<��s�.��^E��S<��_9pM@�S	v��8Rq�ɲp-��ft0�'q(���	m�>�ջG����ܺ��i8���G��}���=3_g���E�\s!3���6?��mɽ8��&�8ؤ*qa�n�
 '�CA��MplL���=Ӿ�y��[
�r�'7�SC�;�v��&��%el��� � ��}ǟ����%�'X���G�%Ƅ�����=�E�Z+M-�A�����,Ș_+�Pݛ{�jt���<�&	\��>~8�Q�������X��,v��4�Bk��L�3I�D^l �\P�L�7�4�Z5���Y�1�-��S�!@w�QR���ג�]�hϼD�7(�Y�bj��gS�i�G��o�v�;W`3���R�J�>MR�7�W
�s�D�����t�䙴u����Esfbb�cދ|�:@TT�xu�@�e���w�����֋oq�Xď�j�}�|��h���_����?�^+ =����0
�����0LŐ��Ix�%�=js�ҫO'y���R�_%�i�h�#�(�$,�^i�V��g��(G�ff=�C���)9�A~��;
]&��6�
���z���$�(��Y�iKk�l���T�DOW�e�}ɨ�*^+�,�̱�@��{(RFVU�%�:}>�)��Qa�L*���θ�rxeK�	�=���%$�@������UZ���^��'�;X{�8��_5c㔅?���^j��$j�@�0�T��+��L�TE�XΡ���[P��	M��JfGi|S�����+�ff�5�tl@9���/5��c�ш�Fe�����^�q�2xD]f��C���G�t`�h��a�q����BU���!�.�j�9�?�\Y�7e��R%���f�cWo��U��|'�+ȕ�O�n��` 8{Wj.,�3}�FI؀�N��J�N)LK��BCQ����U�?Σg��r3ɮ,͆~ՀU�4?�3����m�Z�hO3i����,!d��he\�� RM]�v��@/X��:h�i����J]�D�)�E�	(�d@�~wl�
����`��"ҳ�OK�ɸc�*�]��������:���?�d~ˍ'���f��aNG�K�c��S����M��F\�5�ث����G/�˚�4Oj�XlxVHYEB    674c     5c0?��8q�1ME�:�B�!okjp�X��X��ąV�p��v�Z�B��Q���.z/�eX��w4})�P]w���E�D�>�Êi"���c�+^�qk����}W���Xc*�;A^tHbB^ݛu�����eov�q�6�qU�B�O�+���	��p�`W���T�ލ4��Ԥۦĕ*\��C� {Sș�]�f:�hڀ�cA��H���2v{�B�I&a�i|�.�QH�m�@s�v�8|���N� P�>�ْ�P� �`�3�#�~2K�qm��p7A�х�q\��i�M9#�G_�)(�Z���2���7�s���|'��|�Z�����(Rc��L��2P�n0"��?ݍo@���C�Et
��eo�'�ǔf�P�
lYծ�Ǖ`�e38�5�9����&&�1n�>�7*�~5�D8Cle#���j)	|ig��Բ�飖�G��dQPW
o�W�bn�T��5��O��X�eE���\��ؒi�hh ��v�!�����N��`!T[�r����QB��9r������ٙ��.�	�nW�D[�c��J��t�L���.���6pj�")�����5�p�?�/´���?mq�*��B�/�R�V�u]�&�=
��U+�pd$���b,z1�G@aۈ����e��ȘK��ľ�_cI���̩��C�,S,RC�&�s�����⺮ȗ� �����Gɕ)G_Ce����<�"���v^�����Ÿڳ�?�޴?���e��B=Jt�8`��U�R�X�iXIY����c��Խ��H���ؼx.�A�h����*�z��|�t�V��A����먡zl&̈́�(dh���#tZx�	1� s��M/N���S'w6|vYWϑ�uR$T�Q�!�����^�<�Y�Q��<0i�����pI���P݉vl�.Ѝ�|��7�6L3xL�Ìo���Ȧ)y�̲*hז9�ҡC��Qe���3��/
�\!�#H�MS��r�Y���\�P��j���4T=}+��%d�F��Oz�1<R
�| �J��Y0g�pqW��XD�g]����Uh��Q��/��[�B��6�ə
k_BT���Q��?�
�"���X���[���>�t5�![��ׂ�	�0ӗA\�(���G��
ΰ�+I�<T��J=8�?e$0M�R�ۤ�_Ͱ=�f�fѝ��Q�a���Qs^�k�Dl�T,��f�-�b�n�8υ�^%m�������F��n��D7�4�d�0\)���:M���I:���r����v�����D�veb~:�)@Sr1n��8�ܔ�q�m3փ6�ʠ\�ɟ9�%g������3J7_���Dm�g�,�f��Az@i�r4o�< ��/��*M�v�g��.���:"���B�*w�%4K�;�Q�x��_�?3	�#��ۊqB��Oƙx `��q���j��Yʱ 	ba��PA�PS3j�.,X5�