XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����a#)�gp����P�8����4A�j�VW��vصl��R�PVbHp�&�4f�}�̞0��N%ӸhF�偂����]xy=C�x�����m�_g�@:��|�4����|gA7'�]N%�N���2/��N.�K6���	:�
���L�}�m)�]����V�����_ e���OZ�S�%1��hWez�(f�w[��x��&�8*���^�P��PpJX�l��Uh��9������=�f�������KL�J�UvP%{�E�z��`8K�F3����F5�0�y�j��Xw��7e�
�zܽ�`��HDxlk�	x��'bB�dhUP���<��O�T����G~��F
�d@��1%��{X�6p�^�#�o!~�����c��٫�0x��)��#����3�O��� �P~��U	6D��F���̓dW������60��S�ž!�]��1��p|�M��N�8���l�9������4`)�h��I/�4�2� ��F�I��C�s�}��@r�����	��c1$̪:� '���£�%0\�+,�p�$[D�]�~@n�;�$��a���JQ�*��K����|myp�ϖ���Tyl6Pd�V�ץ�r#+�W@ '/X��Jw�,�W�ZP�+����5V�֒`y�M���H���ąh��ܼ"������̥�Ż?F��G�w�5<�Ή�
+˟�-<���Q1MV�P)��{1�j񧣢��0𖯈��l���l�g�sX��,��XlxVHYEB    aa31    1e40́a�ă�D¾�.����x,�����7��|�]�F^S���B6R2tu���?(��ǫ�;Zzn ah�F�������v��;C�R�������������(c���5c�'n�B�o�lŬm-�@�I���4��˲U���W=�KObPY<�%�3מ��A	- X0i�_�Ni�io�,(կ9fT\���hP|a�7�6�GU�{&�#5�CZ�0曾���� Y.���p4�,��$�v=��W0~�[l>q�����
�l2���j�5_�>�o�g�N�2�J�7g�����J��g��{;7�k,h�B���z47Q�E5� ��~��,��NG�y^��r�&�ޡ�~���3�Z���6yT:ʒ76���J5�JK"*�_�B�-ʏ��c�0�'Mt��v�A��P���U|E��1������'�7�[�\4/8XcF�Q<ٯ8E��+���v��vX��*�&�^�Z�Q�[���?�1�j�۰�Ϻ^9ġ[�
�H�Q��0֋��r�j����������xJ�1��a���}�*���[�.�4,b�9d(�&0)^��ɻ�^����Y�n��:e5��ъ��4K���H��|"��	�Y�K���p���.���	�QQ��ʜh�u��u�I ���K^�����TV�h�K՘�+곷9�>���B�:1&cn}�j�$n�����k,wZz;夌��>������C<�����w ~��������c��Ғ�M��j%vlD�T�y}�/�����"j�.�C2�FN_(֒S,nC�>��Å���,�������]h�$��^�&�)���|�1j�ȀG3%�-�u�oό6��`Ea�cԃ3�(���/<�p��sJb��8H�qI���$�io.{�H�J���c=�2�@��������O7~)�a��+`)�,,WV!�w��~���r����}L���ĶfC���#��|�x(�����h&������Z@��Q���t/��ګ��;�X
�f��X���B�j���)��V_L!~�?W���`Q�w9YE_���tM{�o_�=I�
��4I���p��v{�n2���Z��G/ �r1aQ�[�[�SW7x8q�b�\��������f6������I'E�M��$(�h9�r�A�&E �����/���ŰpK>_爗�Л/t\���N���I�o�}�4�f�5&�ۀ�Z�A�T@1�&0)u�u�~�2�Lm�ZD�����DT��r��ML`G�m��`�jT߇�Vă�Z)��l`c�M�-e�\��qu�
�J¼��q�;�����S�+,e}�/�r�ẻ�&�$SF�LJi#s���P��<���_+�z�Q:F��&l*2c�Q���E01�f4�_'c��s��]Mc5{��i�鐍�RRa�,d�����y�W�dV~���۴I�%̎�8>iW@9��ǯE�6��>� �v�mDpK���A!�׸0s�%�|��VaN>"mf;��0A2�yW�~3�g�~d�1�Fut��R�҂��{�x{
[���uP"�Ua����bEj AT��I|�R�o��8��﩯D%���B�wC�@��Y9Y�jg+;��l��`w��2��b��ϟ�s9�h�y�suSUC z�c{�s%aR���1���-Ӏ>�U̒���{�����Ν�V��4q���5��u�R�7�Ar��*r��p��Q���y��9ϓE�8s����N�"�)7��AI};p AK�A���!�n5��(�q���3����!���X�.��yO�|��ĵ��M��o�D2�Z���5%JL�)��M����}��Ժ�h�x�FA�z}aQo�K�2K�l����o-��љ��F�-�aw8�b�]��~?�^�:*��� ���_�#�J�W����k�11v$`T����`�ӟ��_�:M�U���g��}�� ��n����P�-Z�%>�� �M��A,��eq�"��,�_T�Z��)���6"��_��Z#8�����5�� i?Yo(�ҚVM�p�z���Սo��0�C;�;�_��s�xϕn������fN9Ɖ6��l��}���便6�bĸX�@ y4$nP�Ԃ�J����&��T{\�OTb!�����&W�H�g�M�S��c��A6�6R8d_�6�<���'�{���4�\t���Y<fQ�>$�� �m:�߭��p��r�zT7��u���f�J+xA2S�=k�L�@=�iW�����Ҳ�J�q+S�(
���ޅ�~D@5G�/tDac�U;���6��AGx�����:��7�������JF�K_T�8�����}�V�؏P6�@�ywZL:��'Iu&u5d[��f,Bڽ��yS�Ղ��}g�����\��॒��k�Kդ� ��4���]ŴL���Ec�Ѱ�_�N����z�o�(��s�MdjdojN�9g ll����m��T�K�6��'�@|�EM&l�&)o��x�˪�)M���&ٕGސԟjI a�E�[�?�k������҄k$d�1�Ȗp��~�'�b���U��*�Te>�.10R-���ݮ���xQz(�J��e��*(3��|N����A	TFB��O����vWR���]lYt�8[FH�j�����!gf�,ӗ
��f]��U�c�3���f�D���HM2�3����,�5��y�v^Hf� =�̝��zOA����G��=�^��d��J��kc��ʤةZ&7}�sM�*?�_�'�l�Am��ʄ�,��ɫȦΙS͑Tw���F�(�x��X��M��a���.c_q;�˿���8>�$�$ĉ��=��%�3���Wޟ��ZLx"���:�d�w����e\P1onu�`+=Fy�L&���"S��V���r���͆���\X��;�֒U��2]��h_a�o�Be$JYƠ3;)�Ϩ���W�˶^��%y���NB�+Y�P�J��!�C�t��Z����:U�I��H �O�'�VI�q�Μ�Zy�)���O2@g����G3����/V����SI/�V��0���**���g0�̳̖��\�}2k�Km�n(��[��F�����j�L|���۸��VV�k�ޒ��JH�=�e$��dY"��DkC/�1A9"�F刃d�S�v���C)L���B/ra�Ǎ�Z������C�������gkm������Х��Ԟش2SD�J��rs���La����"���~��w>e�(yL8���B8�X�����n_M3�ޑ�Q48Ј�Eh�}�o5�T&(���r�p��ǿ�D�ϡ:�\�in޸P.���A������)��y�"�qOv��Z-��R��y�B�����ֽU�9��'�Ν	$���{�@���c�/�YQh�l��F,�����mz��-��Z����<ꐹy��Ex�����I���_�t�9�
�Qv*�k�$6O,q�l�9B;ɐI%��
�!Ҫ�����!���PP��+���}���[���-�5���� R�"� ��&4:"2Ǚ�$����`�<d��a��7.i����0m��#*m[% pu��o���˾*�B]�Л��ު:�[x�	iC�n7�M�;6�n�O�+Ⱥ����*�k��s�r�Xh��2�^>�w�Q�~:�}6	�;!�EOF65�L��[4�^T�
��	Ls�p��8�����_z�7Կ����X��mKvcg	�Z}Ԃ�Tw��svS�)Q����2�JnƓQ)����u|��m4v�-�]����)ZN�&��O�0&u�h'����w����l�Vih�.�T^�w���&�BL���,��76\mP��
��	RH::V��V���0�km
ka�fE�<�T��d��	���]���<���0O:�7�~�� ��Hv�~%���
�����C�`67|u΅Txl����3L���gW����2�.0����Nw���O�x���ߝ����5v�r��!��[A�!6R\rZ�b�.��`�;I�Q�2LN���;��o�`�F9���gLY8���i]�P�d�oJV���Q�S��K��mI��R��*�:ޗ�,��18��]���e��-�A�Dς���d�/�C.7�@��mk��a �K9w�$?���
f�7��/5A�@��<�n�.]|wl{V��6.X��������w�'���k�M)w&�X��
Ⱦ�W�+]1�z������V7�Ӌp�����."�/�"�7[����q���_M�"��W�M��hIB��j�l �s�"�i9�b�o$�ϩ������ŋ�$������l��fL�K���&�������s�1T������z�2��cz�H3^�����[�����(���u��2��O�w����=bX�3�5$��aPt�q����D��4�ŏ�鹽���/X��U�
��^�%�i�i�h�Ti���P���T��i�o!���N�i��#�d��Ϩ~e2G��@���{�i|�EY0��1��b"׀�ɯ�U_�����3zU�X�異��	y�=�)	R�o��D�t���t���L����$)`T���ٔ��1cl
"WB<�Eu#��ښ�jD�gjn�ġI�?�9��/wJ�q��d�/��sr���ܽ$,e���L����{���4B��j�x��*<'�c_����ļq~T�,g7N�mB�
{�9˜c�;jn�5E.D��Ox��!�Y���=�0K�a}��u:<ȹ62״�סn�Ώ�z����V$�@F
?�$6#WA�K3zl�ϓ��n.��#Ek?<�Ps.Yw,~�G S���W����D~��f���֧3/���Vg�L.��XW���Ẅ́F����.w�&���'��2��ԫi�Th&i�=,eA���N���=^%i��p�0#�n@7#i�m��;���n�U��xH_�=��i�_Ν�@M�����֠6��Ô.n`;���ҭ5X��0���a�T'�%5�eK =� J���7��f:p��ɘ���$��HmH:���ԩ�^_�d�����?i ��J$_ߓ|0�6�ԭ���������?��0��Z��Z�?��`8�;D������Sn]=�q�T�V?N��xg �w`t0e߅�����[)�|�'	��o�?�������#Z��ɰ�gLYh5�Zƃ�T���R���5� �  B�ҡ#��I|}�;�E�] �¡K�B|<���ՙ�y�"109�ͤ���\E��0;��ax�:��P�G�+\૛�lFY5��&�r[Qo1J�\)%zR"���M�L�w]������V�4��@�}unȌ�hz�^�jt>|uuL���6$�;��"&-ݨ6��j�u�$�j�F:��ƵUY��hRa�K�؈k�k�
�O'eK�� g����v�z�ٿ��$J���s�?#��͟-��~y�ӛ?���%���ડ��~W!�.�!��a��熐�DTd�B�.���y�e�V���dG@��3b��d�&�9��Z�k$W�N��bӘ��G��g¬�{��ы����5�ӽ�rC��k��̊��PZ�S/j�٫`�h���Q������ �a'�V~��0�0e�B�N7W0<���������5x�z��6ޥu�����]:��&A7K�-�c��Njq|@A%)�ύN��6;�ϊ��:Sղ������C2S�0
�Xѕ��<�3�E)���Ek%\��]��c���`[�P��xo�+�����f&�bD� ��~��X�[GίF�`r�T,���H�5��x�����75�Tg��R�,�n��?^�JZ�%�����a��D��UFp�1dG�=�4��QL�ո ����N�6D& �oG���"����Pl7�a��*�o}�Q�����DJ��q���S=�9xN��a�'��� F6B�>���G��qVs�3k���C�Q(SO[��*@�&��t��҂[�ߡ�V��-�5������$����"r��n4���qf*�>�S�+�\�M6�Y*���;iSt!0�y�F�*8v��.�jZ�C�L%�@�7����G���YG�f8thx��JV�$���$������<���Gͣ����W��~4R=��v�#�/�b�.�:Z�gY�n�U�	1f���!�9�.G)t��� nL��E@7t�f�@��qwԡ���xf������b>���^��o��� S��1�3�� 7��MBN%�Sr����#�����8��bk�Ё�څn�d���u�zr���&ܣ�HAQJ��?\ A��L�����������`���&�U����J:~���0������|:��\�F6��blw��儏�j�*�_�������`�ƶs֍u�a?K 1}��%$:���#$UZ��͕����:��Ϝ9V	�rD�{���H_F<��:Ԇq�����7�WTgzy�m��1�ч<���g�d<n�sn��V���������SG���Q=��M�n�#�FPq���7�-�:��YXR̭�> �+.xE��e���G{v�J���E�&-d�^[��ʵk��yUna"�w�8��.ٗ+�~�e��V�ʾ:�k�_�G���.N+���o�EÄ��̂)�e�Y�ǭr�D����j�f��G#m��wxe�'�l�A+�V���B#��ы�b���Cl��`!Q���_�@ݟ�+�it^���n�T�]_p���>*���r���OgP��:+9��G�iy6���/X�����>�7�.���fts�d�c�#E}�,�U�&�n=;�����i^���Qh��S�ouK	�ԉ^=�*�� %s�� �j�V��ϗ�"�*Ժ��u$7�ꓥ{�E��#�W�[����:�ѕ^v�G�O�W���
X�=W^i�IE�b#����yfm��Loy�ݚ|���A��Ŧ����z
`����Y�(*V�CN��Ik����gN�;^Nf8�h�)��>�9j��A)���L�R[�K�>��c���nȑ^�0t\��,� F��M�1�f�FR�=�I��� �y(G���JT��)@v�O�/�@����%O��&��`K���O�1�o�c�	i�gD���ܞ���`��C��g�]H}���y*&W�@�mD���k ��jë�d��m�m���|�/ӉjǷ���Z�ڮn[���'�+��*W��'�Z"��b^&Mj��7��Ю�&�&դҺb�&�+�.�h 1�	��钩���D���[���i/�#w��67"�N �����#���������D&�΁K�rWV��Yl������)ywk��>oW�2��֜�������M���>��bj1��8͆�2��p�V��Y����-VéH�	�6���*�2\�ll��)����jY�#
������Vo��x�y4���<�	����D�YY�S�Π2��o\1����!����ޞ�xB��(���3þ����@d<�M��	�K��;{):;�,"<K�:H@���G9e��3.n!'i2���]'�]�j�.��N(�n졙�A��q4���@�\��MP�{�ܔƙ�DF���q=�-���l�0NR������Xfg��f\k�z�7_���;�ը)�CƁ<���!˭�NA��=�8+�V�#�}��*��$