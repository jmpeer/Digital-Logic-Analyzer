XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��G$�X�xo�������B3 :1��ŕMo&1���"����(ʟyϬ0�Sn����w�8 $�6eB�M�6�L�3�I,���t��)>�-�`=W{:��R���oB�4��(2^��\���y�^�բ/�<!H���l��E�9hrlt������@�`��p�|�l&�C>��ɜG!�ɜϗO
9B���o�_��fL�_�������5Xހ��͚o�=`�aJv��n��7��{e!�lӇ�=D�YbuL4U�^cUJ�(���A�L��k��
�fu�Ink�	T�=z�����}g7���^dx?����R�u��v<���� �xx���D�ɰ�7�� �X����JՓ�����L�r�`+$��>4�������+XJ���;� ��~sɽ׫�R�.H�9<��ʏ4�E��ۤ�C9~��6n�u����������ؽ�#�F��?f?M�T~��2�k
@�J��1t���&�U+���Ae9�=r�-��@h�0��x����J��Y��<�&50s����y��w��e%�"�H�7���e�u��D��|��-����G@Tw\��}��M6r����d$���TT�ݫXN`���~#F��#p��KDǚi�CA~�����ek0n�I��^N�����x>:�9Oi��aH�ӫi�wH�=7��-|mOK�Q*r�3��+3	�zum,V��y�eTK�ݗK�ܰ�2����˚,n�4�?�P����c-�ΥX��9��B��\��5�XlxVHYEB    aa52    13d0��$����+#�ӣM��2�ѹ�����;���T^��{l�n������30�eΛ7YOE�~,n�h�88��F^c������"-�:�������s�s��rD�!u˚|�C�<.�ռ�~�R�S>�ÌR>�/���n����G2�,ƨ1��Fddd~���)�X���9��/9O5�xO�ҟ�*��{+{%�(.~��;q}��������WfO\7<H#E�6���Hr-,�d��Y�5����hX�E?y:g�y�M���m�k �Bmv���]g,x��]�()z��$��p��|wf��wq7�&lz�u�k]V�v�Zy���G9�1'��eE��7g����v_�r��M���x~�1�[\�L���M%��R� b\Pa�dlXA�O��x\���ձ�G�Lb��ɬ�`i�ِ:�A�NPӭϥ y���gڢ���Ȓi�y�Ӹf�� ������c7odI�\)��i�r�U����Z!ɂ,���v�B���IIX�`p��\��z5J�u�jBDnq��v�K.NG�6.���X�Y�)�%r���j���2���'�Q�%�PPh4���	_Ώ�3�b8KKjgﵩ{:
�L|���D�G��/?��D�o	��C���4yդ��9{9`�m�I�B=-�F���m�en�Jrp}�k���� ΢�7�Ш� ׳Y!�z|�Yn =3�� ��0E\>�$��a���^%���1���򀰍ep���n &�I7��17�����#�<B�"ъ�˺���=sY3Q��!����F^��S�<o���Ǎ}`\��1~╸t�a�����
oZ�ȗQt�f!��|�M�0J���_�v��Kv¨:͙.n�4'�w�+�c_=��wU�Z�U ���fO����l`�'��9P�����谣�!�.8�1���;�X�Ѽ����������.7@�13s"�����C.�o<����[���f�J���'>><Iq��C�i#!ۄ-G��H�G�׊�qBt���AW���s[�Y\���+��q�,ը���B
p4nޗzP��Ch鼐��RI���<75��uֱyjTG+-�`��Lck�̯�9�\,�+��W��yX��{�I��?���H)n��Pry�@U��+�ɂ}Hs^����+��� N�	�$�̓�F 90y�t@�,��!�_�%.�������'R�7�=F�cQ�H��LV�"?�~c��L Ɛ�s�Q��.����Ý���	4+�F.� m�9��󆗘�ڟ��$�)8@�{��ӧ�_C�*E����n8�����)��
RY�ew�� V�qi��$�9AQ���P9��.�)����=;R���AS%B��@�n�U���X�6����U��-���a�����g�� �N�- ���w�d6��L3�`�˹��#_z�|1{��U֧)]���@m2�(�j��>_�\�� k�_Y�e<dOP ���@D��QK�2SV�I�ϋ�{���R�1���e��Uó[���1��^,�B�i�}�a�
͸��i��߂`�����$(\�^+�3|z��.}�g4���Ҏ!��7�ğ;��c�1%�E[�7CS=��<����v���n�[|��� �ݴ^�ix��C�Csð�"\�N�Ʌ�D���8���ji*n
�)n�J�|Hfjz�Z4� P��n��K�q�q��E��W�5�	��EӬqL�����B���h��q67w��#�AU\CX� {��ܻ�\��]
��`�]W�>��\(:����&���!n��j<7���[x0
��:V6�x�q�TB
�<�׾��C�E3����"�PL=���@uZΰF�Y\~*�(�d��:�U�I�"�V��^�C���5�_&�X�4(�)��ж�&m|O�����/�Gԟ�����r��|8�h���E(��֑5Z���_	g���fb�/'�ϝ�	�S}L�t���/��]�=~й�	P?�%�TBNY��Y����aAV���y7z� ׾�Ar�ik�|*��%�Q5Eo�;:!���S��?NnI�L����5Z��dBS[�R9]��-ȚR�)��J�y�3���-,�a8y/�ɘ�K�n;o<���;����-`=�y���)�ts擫7��둱����=��V�}�M��/ ��n/�NX��bp�_�I1���?�SvT0t��<���vCǠ�Ϝw �=�P�V	Jl��>�
����~>_p���#��|n__��?���x��4]z�n3�������:^�iI �z���-�\Y�����|P���YyPutn��g�(�xˉ5sO@C��[�/�}T�Dk����7K�8]T��&9�T��@�릇l����--e�ڽ�4��5!TeB�W����n�ĉ\��:�w1F�:���ipׅlQ�]����B�c"<Q8g6Z�m�/�v�X�}��ɇ�-;3�k�$�9yB�����t��F�.|D�)�aR;ڋ�V1{�T�Z�J���g����K��,���)� ���)��lz�5F�����d���|CFV�&� <�D�$ Gnl������,�)�3����� .�5x
E'+~[���$tV ��*ͬ�+}��g�1PX&� ١��E��՛���nd�	�v�BR�,���r�s��WO��U}+�$�b�����$�EX ��[z��_�K�56�s���^J����?��B�f^�JBn(�p���[3�:�(X#�JŜO];ӕ-����!]��#V�]�Sx��vs&�&ə_��79f��Η���z�� XB'b��ϻ����X��
I1RH�xL.�Fp�Z�>��J6�_d�7��z?�f��Cs��9�u�_�����4��c�7�gl��_��1C5�M��?B� 9a`e*P{L�F..e�������&!�۲!OY_������9Ԍm�T#�Z!<-�T�#�tR�+�^ZDꗻ�c�{=��bNT|���D��ӕ:[������w\�9�1�=s��Tݤ)���!�@r���x��2�6���:Bv0<���5�$���@|И_@KB�3��a����L8�.�$�oP?h����t�G��q��59Y3�~tZY#u�� Չ�W��v�]F��H�|�b
j�iAܑ��>f�G^����\Wa@�?콨?��
�ڟ��Y�ԇ
-թ��
	*�،��/�� ����G=E�O��`?�ܖ���%�ȱɤ�%g~�&6��۱u�"���(ْ+�8J�8�;6����Wv3�]%�9���`�`�-��
�n;�R�=��Ht��ɋ����BU�����rT��7PS�y�n��d��$����X���}8*�f��P���������κ�f�?��Ö���Q6Xs}5F��y`���� EF8�$�H%��N�5�KJmY���p�ƙ�3��P����N����&�2mՏ����"�H��ieW�Le��D�[�Y�?��]�������G耣@<Ȱ�fj���w�U�ٶ���p��d�5,�:7��n�Y8F�P�0�X<�:�Zh�Ԛ�R�h;�(��b�r��\2��w0�����Pn�ӊJ�K�X��1M�'	(?�@�~��/�I+�R�Δ��Ŧ V5�5 �Y�=���r��~�w@��mB���}��$*��1���d�3&���o�-�����hz�Aoy�ED��A=蹦!�'`��o�}��J�	.��Ԟ�����Wϕߤ�q�U?]�c����ψ][��PK�]�6�S���|v�s � ����OP����K����BN��I��н��ϫ�����4���9���F^���-�-���Q�U_}};��1ir6!����Y�������ݞA���u'A�0U9����ؙ���q?㛮j=�<ƔF���#�zHG$�A��f ��G���]7&̢s'}ؙ2�(q*M�ƼLJ�x��>HW�u�%͜�k��Z2;;�z��~���`�#���kOA_G�qZ������u�*5�������\�.�+���l|?��'�P�>tc>�} ��za��s�a[ʈ�Y�3
�����\5H���=e�g����2_����6I,jp�8�0|����aƧq-�I�������(-��=�S ���pۓa�6)խ�U�](3Дd�'ᢄd�+���:b��R�*p͙q^l�	m=�<�D�v�TE-�x#Ql(�4"�^6W�$��pL~ץT/Mt�o\��i�sP�3�+	$�nYL1�,�Uy�	��\uՋ�Y�l�u?FZ�i�g�(=�TXGq)����=��� q���ҁ����]� j���eO��o2B�4���6':##d�ي8�b��{M��
�>浱�����Ը��1*Bz�2��ɡ�^�f�Tv$� U�/�`;|u:j�4Ʋ*r�ѱ�B	�b����^ҏ<���Kp��QD`pH��V�1M}}gm��0�]��1��d�=��_+��g�KU��p�4#1�h�PVS���ϻ�պ�,N��(�����y�0��U�C���haa��9W���m�s�l>� �$�)�� %���9��o�y��LD��
k�ت����l���Gy�2|�L$}�A�0D[­,��M��e����6�ʓ�&m�xӎh,�:#E˳�
`���	�5=�SRз*m�+�|d�E.S�����fQ��CQ��6 `T��Չnq�;��̚ /���LR���<�!�B�ܢ�V[��~.��@z��6_��"AU�H߸��k�%���ްv���pK������|(�.�������/�T]cr&z:Y[�|���޺NL�BD�++0la�#�r��T��rI��g��A�Xj��E�+��<��p�U� �A|Z�S�b96��}ī�	?.� "͍aG˩u����A6'  ����H勜n�=}��heÓ5�i�4�F!�n�:@���[xo�a��F|