XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����^
=�2���V���H
$Z3%^�6�h5��k���6z6?���/]�@%Z�Ԓ��;���
��b�����k�#^�8�<!1�U:b8�CS�p�t���N�V�f��C��tI-��X�ɼ#?��s�f�ڨֆF�`o�f G��ngR���";5$����ƑS���JI�΁zFŪ�l=n�f\���:0�a�$l`׀0��w�q���*&��91�h}5��)�
^W��!��A�`b1]8�+�_��?Cb�BY����r��d��4ބ�9}y&A���� &�|��I�ڶYթ$�}��j5X5��p=�J����%������L^�d�]j��{-�݌�bI%�fb���Tt䷗95#�+9��I$�p���w����~�ޱ�7z���M<8��N��Zt���y���t%��g�=��9�%/@f̻�BX"t�Xg �)�ըY> ��")���}�����޼�|��P��4Ս509yI�`f�uPaӹ�d�%���2�!zk��tt���V2������)��J�@Ll�=�TA��h�oJ��[˔�h��o ��ؙ�\��
�b��|����\���L�"e3ʣA?�ߪÅ�"z�	K=�6&��d�K�n��U!�Αճ-BsDe��R�͔hd�_���i{bjM6e"Зw��x��m�XB������|2�4V�u�m��p{�)�#�)|�ZF\����i�[�ڊ^�DG� ��?�E��l�<xv��)AXlxVHYEB    fa00    1fd0V@5ʯ�B<;ʍ/�.�J+Z�����JRK��EN�����=k�G�d�m� �?2d
��<r��ø�<b�(Z�(Ƥ�B�-n�hG���#����"i�k<٬�[����.�N���ծ��ޗ�|1)0����p�}qQ�6!5UzH<����4�(�~*!�`e�m���u�^���i�b��&�|4��!�!c0��H�X+��=zCXŉ�����P�4��4���tW�9�-�%�C������{?�USD(t��d�.?�XM� R{RN�8���1fltl���v�Ю����%+���d���ʅ�(m��o���Y���N��tk`R򂼲�˅�@ �ߘ��?;*(��x�g�cbc_*��d�:�Ѯ�撠����e� C�={`�S	���������5(��#,2�9K�t�k��B1B�j���M�
�����;d��W^��U�;\�9n���%����42j��ҹ̮[�%�$K}H@eSPV?������t��p��B��"`t��p��g�3�����K�ߓ�mR����%pT톣�\�\I�u;=0�MF^O繖��gCQ�Ф�(/"T�p��j,��P��s���O�cI��uL�#��
)r`��C¯���㙴���5 �꺣D,��o�a�-b��V�t��	�}��'vow>��ƴ]wH�S�Y�t��>�;<�к%'�۬���#) :>�{+p��=8�]�Y�ܢW�~��]HY�+�%��.[�PMŮq'�<�Z��u�M/\ �Jc�w�)RT�1+�Ja���@�w��������~�[�,h���rG��߾�L��)����x'bQ�f}X�#�sXD�L�rQ8x���Ϙ���#x�c����;��fuV�Z?��!2�C�XЂ�T?.�lǊ�{zD���r%eQL��QF�Ys"�|��ZW��^�\,��_�}/#�DtP=�^Ϗ���ު��ʑ��h�<n�%��f�������BySԞg�ѫ��,�� q�8D�BN�*ؠ�wu�����Qס&�D�e��-^���ո6Q�AV4�f��ΐg�P1�t��D���U��M���e�^�+]�����<5�_JN6�z㦚�`�����u���2h��myE�C4̫봾�.�z���:����..��+2�
�̮6�:��G�b%�P���>i���Ir��n0��K�ɎnB�o�3���� �r���yyȗ�r"N�+<���=Z,�|T�C|C���)B�;��D�֑$¦��v��=L�8+�.�:m������[D��.�*$�ʉ�ʣ<H�8��Pgwx�����^�є�~�+PT"���W;$�󾛮�f�0����S�{�J��d��hSj4߈��dO6~D%�����ug]�B������
6�Q�^��cTu�|?-�3�1WPd<���˟��Lؑ�Yj՞$JAK��6�LJ�R�-�����g���g�9��ۋ,��
&�:����E2[b��SQ�~$�Y����9�
������o���\��0�&C�A���-b
��+*Z�,�g������m����ڇ��>)>U��T��|,v�a`� [���c����Py,>����f��lW0Η��h8	���ƙv^�k�ha�����d��AlW�4`4
��j�Tz��y()�$�qr�A �3����k�I�xvB%���9$38�=��)������>�V�~���l8����sr�Ύ�s7$��N�}�[�{�h�`���R���9G8{%J,�N��߫��t���2��V�Vi;M���g�.��='QP|��=^8l����ŀ������Q�Z��:E�62��g�C'���'yU=���wGĦ��$�']�}m�8�:�HL'�|��ɋ��V������l=�۹Ց$5��i��� yw�5C����\/vj��Ц�4�9~� E�fx:%�m�t�gw�nd����x�;�	���Ҁ�P��k��<n��n����7�Q9_�B]��d����~1H����M�[@U x}���>��q(���ᡘ[ifø�P���T5��OɓbP��S_Ff�g��>�쟍>��4��9�(���r.�+.x�{�A�g9~4\���hh$�-a�A��?6���3[x��1�x�UU?��Ўϛa�5�i�-��g�
����t�U�jߦ��G���U:�1�c��ǡ��4����s��.��r�KSB��2�f���IȺ���i��BN�Un� �he%��W��.���� 前q���;NS4�?hW�	��7�vhy��#6ٟ��L������m��LN�v{��L���h�#�]�t�/�+��i-�HS�k��N����&�2�嘿$x@}��k���M�Xӵk�v6f|�P�����L�۩c!�n�{�YR)�T�cs2e�2�4iK�җH�{�wZ'�b��t-��޶���������Wk�<���S4���/H4�:��g���g��=�_�Ƙ�#�K(�������t�ш������`s�y���(ŽcQ��p|������U�?��d�Y�E��]�Ċ뻢�?j�ڧ���2W�����+���rvu�y��՟�T{���š��jcsyBt��߆��/��0icܑC�'>�����z��<��$����\�{�xtD����`����MRJ8����3����q���AK��#&��3��{xu�Qvѓ�/��"�tc�t�Chdӎ<W���}NRޔ���@��'DS:BB�y`���z�ɝ�)��B�)|$��ww��}�7(5��*Y���2��4 8�����C&rU�zR5�T�0���|������=nOB��@���}Uڞ_�9x���dNz	C��|3S�X��uM�`��ʒ�O��|�l��~�eڰ��{�������_��͆b���Fk�ê��E{A@�-qU���%�rAL;��N���q�2{X;_q���4�E�9F�������%����Ӯ9no[_QǄi2����֣* 4I��ܴ1����"����0�"�|.��y��$�� �Z��HtL[��A�L��b"4چҏ�zC�*��������g�Ո��M�6�x�RS�����1�����(�[�	�IH� X�XUBE��_o
�yk�tP��ڰ!���a��k��U�^>����ZF� ���q��������%��o�7#��<r��b�u"ObA��M�ˍ�@���V�uF���LS�v����E��Է���w���
����*]��q_m���tLrH�B�B��!Lq�B&���9 v���4	��®�BE��"�ޯg!ʐ�S�ۋ��~X��k��:RoÇ������\���2�)T��~`?�?��i,������By<	�U�X|���N(�H{��S�NݠG��]�e�q�#sc���dz�A�_�o�&7��M'h�/ �maFi��}�^��O�8�F�I�\��*�oJո��[�g�����R�I��]\���(m����A�C7�&r�߆?~�a�j	�I|���u�OY�<�%GD5�f�d.�p!�L')�sV� d0�e�
l9x���v�-�G�UJ��X�!0x�NwrO�A^��n(Rn\�0"�m��.���~�]��˩"�YqY�)�7�>�E>��X�g��}-^���>B�$���F��%���|���!W��3Udn���K��D����Q�s��F��q�Rl|�-9��Z�X�]ĦJJ��٫b��i��nl�4{�v\�J����Ai2V��	��8	u� �)-�?7��IL�p��>�Doۑ�2�x(�S�B�B �)NQ���b���d9@�u��E��
`��(	~���v�~be�w�����M��%�M-/ek�[��{��h����UC�l�B*��m����
��:yIDVeyG^e��<$
�&����-'�.@�r�=��÷�$�Za�	�ZWs%��qI�>����FT�W��V�?DB�No&O�� |R+5j�;+����"A:�ig�V�_!�q�;�D��yb�J^^&A��H��	��1�����Ȃ��Ĺyw�#�/2���L��G��r���D�@�ez2�����F�8��F2�vP�!t�W`G���Y������6�g!���ӐD?^�ƶ�W?=Hy+j�hgZ��]�q�#n�hN��4Ӥƃ���C�,
(��lZ��0`��w͝�,0���j��=Υn?ܠ�w�\��#P�%�M���C�Xnۤ���#�I��L���/����/^�M�!ؒ<�{���#Pq�r�=$s�A��2� �ĦJb���MuL�k�=�u"�r�iz'l�6I����<��G���Øoݳ�24Hsi�pF>���3 �H��+TZ=]���R�Ri��X��R]�s�Έ����m���z�4�H�j}w��m��ګ����8�bه�=:[@��	_�h(3'���/�}?�[%�a!���D9ޝ
l���r+��RUT�A$�$(��8,Ć�n[Kޥft��ς�f�Ccj��ɽ��H��'������Vd�>Hyjp=Ɨ�J��>/����h��~@#��3�'�+R��������5��x�Py<</K:.�VN�5\v����n9VWA�>�K]����|(��+!� �3�"u�8�۞�7. B_?�f_ʧ�xg��D�ٚXP�}	t�e8�A��A��M�4��f�����%��E�$gYbȲ��?������\�3=r��
�ݭO�tʚ��h�#,��8���C��i�j �.T6���F�aƞ�|]����m�왝?1�"sZbK�4�R�����ۃ[����6̈́��A��cqēJ��-�gBjc%�]Q�iI^����!@���_�a
�e�9�����̓�s�ś>d��V :BlQ��=(5c��´��\������n����I+f�ቯ���)�Z����A
2[�y"5[�:��/y�s��T)��qe�&P��ݚ�)e���r��l.k4��7yg����`�k�a5=4`G��õ���;�Q�E��ao�-B�S8_J  �(���6Jf�Q��L���K�SOu��eNj�ti�{�<q��F)D�G�Y�{�S�H);��|= q��7�*���$�>�����Kj������_��;�NhQ`�D�����B�xpbW"J=�t(�q�؀3(Ҍ��iE���M���Z̚�~�ᖰg��Ii@'8m*������&� [�_�H}���ȉ}GP���R�0�.��au�zED��q>��b����'!k5(l�iE;B��� ��2�0�t:cg�J����O�*F�d��A6���kKc-m	�kZ�������I��p�c��*�P��uP�r�M!���_ ���n���V�.t�
ݢ��܉�<!���p�v�Ŧ\sL�!�VC�I�H�xתL_�R Ix�`�p�FΩϦȂ���L%��)��2�&�rL���:b8�#��I�zT�Jh%�8��u!��Wx�'����N���'�ѰN1@�֯���twU�.^�g`}�#p�����36.���\����\J�:�h�J��
"�4.�+�w*��P�&�r�0���ًU�\� ��*�p�WՂH�'�_��%��G�3�K{`8b��-�G�W)��1C�� =���hb�f�Q��qp�K7tI��K	��2ׂ���C�i��O����wYX[~�H@:�s���CD�@i*C����sED�bGoAP4���TQ��� �]TH�׸�[�K~<�����h���K=�kї��w�S�Q�I�E߼�w�4"�_
砨U���j禙��Q�_�2��C6e�D�@Z0�j�{��D���3Gu��>K7ÿ�T�S�ۗ���'��d=��'4��	VEFS.\���6��w$�N!((����]��d(	Y��t
��5s�O!E��kJ���JX)6��H�Y�n���.��ꭅ���Z�"��}��lo�%�z�"Y'�t��WWq����3@P��`�0����o�;s[�^�� ΕD�t�[�q'f7;�&�EM�"u/N�����My�e��
s�n�l��-R\3���&a��	�u�l�x��?�JGB���}��2"��VI��鶸8^UXu��N�F�Ш��6d��Nx���R]���8l�"�y���_��؋�R0���C<��kBF{����Fȱ�\$�D�Ϸ6p�h���."����Q��ѐ��5c��]Q�!2>m�ˑ����G��B��de��mt3k�RB�şw�aW��u��G#v��9���a<�<	������[ 57d�	�B}�}q{�
��^��ڞ��&a�^���m����ם�kGҵ�h�E5��"�:�7���<Ζ���%@�'u�]/�sܙ�ٶ��Z2�v���}RrB� �W������}^��}Lͧ��<Xu8_Ί��١��y����:o\�^ƶ�q?�=��f?���-����='��YEtnlr
Q'�Hq!L�T��&;��g�K{���L��"�����s8��e�.��K�a�a]U���<(\H������7�t��7ݺЫ�������Gd	��tz���r\?�R��콎n1���/���5���!v7	���n�Y� ��]�}q��)S(��� @-�t��SV��?4n�@��~�Py3��ۺ����d���p!{�
E=����A2�VISi�u���$����Ҥj��@�$&ɟ*�W�y��V�g!@=��3��5�"61'4�'��](k����h�F�wey"����d��L� π	/�s(r�n��$ �K�ﲔ�V�4�`�M6�x����%�v�#Ac=.yԃK�r���8]\�� ԗ���5$��T�ֺ=X��ds�Q��$�	���y�3�kց�j����=9qԖ�-d�ʅ�&���;`��'a��aŷ_����j�@=@��x<M�_\���8�'�.~�)M��y�yu?���,z����+�k��G?�۱���t�6gVr�o���i�ŗ/:�TYإPV�s���smeSG[�>���n5|��\*��h=��=���-N�Q�Y��l�C��t"$_3!�-��=�g�Y�/��`�v_BZ�Rh��K4J�a�䆑]��g<@o&��w�)�!ǰ�6�L�"|i���{)��L�38�
(��؎|WY1w�X2S��E��0,�Y&��߭�:�[
�1|�Q�vo%b;��`�dE�8�#W"S�je*��6%mM6Lv*;�@e�\�.m)���z������n�{�d����C���@<)�D5�����{%�m�Dgy�G�ň���lsr�[&v�Dl�ߩ#3���zxqK	ؘ��|t���?�C2�)���<�h���RA���\֌�)�6z�|(�����s�O+\݊Ъl~���Ȼw�p	�\��/��RY;)״奡V<\��T쾖���E�NĊx� ��$��K�8*P1<f����m�*��je|EV�R�bF �q�n�SqcW�u��@q�����F��H�����v�{�p��V:�D�ǀ�j���
4s�f�/W �����1���sU:�ː��1t���>/�z�CeD��/��7V"��t ��(�PA������Ck���BR۶�;��G��T�d%"1���Bܹ|?v��%g�+��@�Ć���^low�ߛ탷��/�L�0_?��R�> Q��Yʇ�<gm&�+<ހ�'��o�& ���#�i�bס���H�NqKd�]����&�}Xj<�ST��6�X1ΰ���sҹ�B�и�!��Q_��9ϐ����gE<��BWE� �#�3m���2i^�LT��$�-����徉\�v��m�~�u.Y��
�~Y�{8i����w�Ԭ]�S)�1U�7��G�J�D�"���Ji�����֍��OJ�Xx���=�ϒ_<��/�v]�Z���S5�^x��0�7 ��8��4��[��Ta��6�ZlrA-O��*�:_$��F�՗<�R-��XlxVHYEB    fa00    1340??�q�k���/��3�h���;�5�������� �� ��.W�&���z:����Œ�툅]�!0
NRgq�8���� ����G֥��?�[f�&�>�F]�-?����*O����"��V��9+�r� ��˽ۗ�Z���E�|�sUNN(�l��O�>W=�6Ѯ�٭ǫyG3ϛH�he��F�Vߋ��I��\��^/���xn�7w�P�˲�*�$��q�����e��d� kϠ�;�B��2���Ms/�d�;��2v��i�t�����d�o�в�	�#4�C���h/-����gR�M!2�ŧ˃9&����)�#�정�o�2�*M�z>�~����<����d�(��ńX�)nJ��>��Ѷ�(Uڳg�eb�XVC�?�	�h4ժ۠���YB�Ka�A��;{�!E@�߉���rS�`��k�s��a�4�e��e�1w2�'�%ݜ��A_㐶�0�u��s���%�|"�xz�GA��z"|�BٶG�(���0�H}�2�k�|��_�5�e�������i�M���(�DS����z�¦ll)������о�A��}��C�I�#Mr���h6�V��?�Q�U_{	s�)�'^���f��X]!�+�q�������G�4<RJ"���	�V  �y2�e�(T����0��t^��9)��6Ɖ״A�� �=�?��vU�^[�PS2�,�9@�^���f���ޢ0f��c}�M�庐T�z(�b#�ϥ���l�$?��ځ	��h΀�*YƵ0������#"�%�݅�e�.�qE������$��y<nj���������V������2�R֨�?/��8���X�M��)6�!90����撆f.�)�c��}��ۄ�xk�,�@��o�^�"�:r����Jқ~J�G�{+�E�#L���*��e�%���JOR�HҲFSr���	6bN�ٿR�>۰��u<R�&�Ѭ�/���'#�ՖB�J�s��+��e[��e���Q!q�ͬ6�=liW�Ȓi�C�j|I��NCqW~kD��������|6�m�Ê.>����Ț���5�7�gD������#X�\�P{�$2�##�@4�K�� 9\�(}�AjS�	!��g�mXD�(���nu�I	��Br���P����g>N�v��Prz�J8����dS���|ja��^O}����t(2.��0��dZ���Nkx��_�|�OW�&����7�����ɇ��fC-݌�ܧe�S���Ά9o�#�d�q�%P�|�s�����4����A�f�0���$btm#�����"�s�ʽ'�,�������9e/�lξ_-��`RZ�2g�1Rr�%dq�=�1B�J/{#��W�ls��fAy���1�1�~O��׮Z�fZ�X�\��צ<4�;j���P���O�}_��H9"��޼ X(ű֙��4~�F
XlAD���k�U�U��V�������v���+����F��_1��t����̬(Ig#��ȜO�E;�W�܇�f��Iܸz�J�*���3��*]	0l�0eOQ�[�;��/��=��� �'�l$k��R`4����(�w~���.Ϲ�m0LJu��9�$�9�6�i��`��v� �s�"2����>恑�j���5%�����'�]-�+Y��r+�������4���+����u����=p)M�$}q���:F��	������d�q�
z����h�\
�����kb_��+�3"����Zˀ@�n%�*g��s��?��ma��"��+�d�)�Cp�II�v���aI��p�~y���f�X�J������W�3�G�H}и�'x����5�<�]K�D��:�@98o����|�����q}	��So+��e��84�����~�9��+�D�	��*�M�}��N-o��°����� H������QYH0���ʥ� ���f�6(���7�|�߸ A��9^������׫&9���R8�@�eQ3��L�"���꩔Ew2ea��,6%�F�`BCf����A���f�Ӡ�g
��u�}g$~�� �3���!0P�D��5�U��P�䘑�F�J,�������@�tܘJ��Hc����{��4����S��>2�-ק���D�K���ʙ��%�5u�gO��n9EA���QU/6{��l��[��¡�;
�'� ˩-i}a`�n罤�"����a�,���yT1�}c�� &���͂m��j�ǩR����_�/ls����`<=*/����W�;;�z^��}\J��y4�
k��!�l���m������CgXb�!5ȔH��!t �bW��A���.X�٩_I�N��{H^)<��{�o�Ǉ�N+[��Q!3wBQ[����X���z
]f%/��ݔo|Á��"���aP�*�˪�PA@����D�7���������2"<i7���Uښj��jD��?���l͌zl8\����K�ez�,�!+��Vƭ�+�t8`��V)X(-��ks�`��}[��a���i�H�7�P�y�iؿ�gY\>Z9�H|#�f^Bڝ2E�O�YU�P�⓳�=' �^�

!�隕W���6�iq��<>/u�Yч�O�t�y <`�*�-�l���n�Y�f@������CC�t.n\ϵ����yN�Kl/m�yrZn~L#��>#�{Uŭ֢����k�K��sE��8&���%[6j���g���6���}����=y;͜;Z��ѐ���l���H3�#
�Qo�V��:�y��K��JF��r��R�XI麁�R�i���g�,�-���uӧ�2�.V.�Ux�NH'I0;�Z���*s�,<J2-כ��_�~i����N(x�ո�BO�$�ۧ����� ���}z	�Me�U�L9���1!˥���0�)+��Oe��=�0%���r���Km7�Z�1MRv�i�ϞB��n��&B	 �����`�-������=lv��rY	2���҆1_����ͅ�d��V�%���n�.���� w�ԛ����i��#q�ζ�^�rf���=f�}~��8;�r�l��R :V�>���D�A�Br((ܳ��ϗ��,��}� �v�W�բ�-f�Ŕ0���!rrѧ�^r3�֝��v_�ESF���ʆ���@���-�?����%�t��b�A������炗/��K���L�T�y$�x��,�`�?x�v���*�={2���2߈�UVc�':���t�\7c42��=���{��`����0DBT赆|Gt���u�$��0<�8j�A����� )�IlC�̫	ye2 �ɀ{T`yl�� �k�WW��^�R��?.�1)���{�z�����3��y�(f���(��V�eÀ=>�.r�-b�A2�(���s�I\cςǶ쵌�;HD����$;��O����ܶ���oDc����<��IL4�.P\ F�><^#� O�Ln�:��T�Ș�/�������^�'j+b8��S�4p�q�G�T��Ͽ`zἈK-����ŏ�u��[0�vN��A���rƎ��ϫ��N:�}��x������u(�.i	GC�N���#8����SIz�D��׫��8���UF��{Q��=≊��2�M����@p?��;+�ߧcuYl�1|6g�iX\��F6b
i��O{�Y�^���t���5�&�;D��p@�rZ�'=���r^��[Ĳ���Zj5᱁��r�M)�/�H�%�U���͊��FGO�l_��>�t������n� 0�@-Ę,�-3�>��·���l���:�%�Hp��Z�6���we�έ��O���1*���
r�4ۂ
�K�!2f�n�LP�Q�?�d�]o��9��Q!b��EL@~y�mhL_��x���M��͜�(q%F*��7��%�w�q���_�Z:�<އ��n֕s���Zi]�C�� ��a�YPSف5/Mz\�Ů��=��Z���kL� ���,��9Y����/����Y�U,z"W�\g )����e�pƧ�bɚc�!r$�,����%}r8~����ㄯ��Nm2��p���E�6�{d�Ж����(��}�8)W�g��j'VZ�v�l�ݬ�5i���A���>�&H���f���ma4����o�L��R���QI�N�����O3�z�O����X@��"gt�__�	�LT\��1��"�/(���9��T鎗�׳A�ꆹ3D���z�� �!i�J�9ۮevp���� �y�x�2̀� �,�:��3�&�V��Ϧ�u�GY��& ��iȴn+C=I*��.k��+@������q�xч}؏t��P��/Z?�nZ����CF���6ob6e3<'��L^�M�GX!�6�� ������O���"���fM�1YR'�h̊.�[�5�$~~�驝�y��<=�����4���5�X���-��ݐ�0�O�e�`�
`�Ly{�W��A�|9ԇ�iۉ���禨�'�!�{X�q���oP6L'=�������P�?�F�i��?~.�N���3G�ŚG\����]����g�K~�5��/�C?���p;\i����1H���iΉ̩����@P��'G���x�͓�g���=�~���;Ÿe���+�Q7��������d�Bp\ƸVQ��˔Db?j���R���������PI�`�=нbs=!�P�74P���)���"�A�eG�zb��zeH�GF��~����ڈ�C^���Д ��?�b���Y�-R	�k����À��L�����T9� �5��9��N���{	�a��꧛Y�cq7��	�����|˃܍�a���h����%]���z�Z��q��o8����g���j<�ƭ�ip���QÑYO{���,\�2�mx,�	�A�1�ߎ:0�a���XlxVHYEB      e7      a0D�d�H�z���${����d@(�;��pp}���J�D��T�V�8H����r��#��@[�?|c�Z�a�V=-k�������ʽ�UE��ݘʥ�O�J�����!����D){�)�ٲ���/ ��'T��nPfQ`ӀkOo#Y1