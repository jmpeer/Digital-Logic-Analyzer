XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���"��->�k�F�C�}gb��R^ w�|)�������&i��mG������4v�3�4t,j�.Ֆ�s���;C�@�'�{�t�_�H*H|&zt��Y��
IS�㣳�M��e��6�&Qa��SN4��a3Kث}q��%`v'i�ٱ�`E�
9=ײ��w��(����-͚cq'|b^U}�����l��I�L ҅{հ�h�sH�J��e�W%F1k5�Ũq4%�c��CzH��=�F����.�����s�X���X� B ���,>�������ɦ�=F�;��1�E�zw��\M��aY��-I�}�IE��_aK�1�"�/�D�ۘ���s!���$����A�珌J�h�äo���}w"M��'�첫%���Щ�t�I������&_����K��ž�_R��m(����u��57�t�-24�x�Er��n�c���\��!|x���-��Z�Uֵ��*u8�K��)�)�K�=��y����w�X"�{� _���-DS�ON5Vlʸ�5�\Hِ�b�����g��f�We����_N�	�{���C�e�Q�^6�ƏǋMk6�-����t��ݩM�����ڟ���x��g]�ʻ3菉;G*�^���!���{�M�����}z�V�鉊��Y��u��:��潟�D��kD�f�on%��A.�3G�P0�)��0Ҁp'0�bY�p�AG�I�A��j�����z\�ׄ�g�НC\6��uNN�XlxVHYEB    ea93    1880�(�ޛ�����H�>���Q��V�0i�9f�4K��[Z���� �5��s&"X59���.v��ËarbF`A�[$�/���=�3�K�T�V����C�z��,���m��+jO~f��0ՙ�����4�n�������5wb�9����Cb����,���t�q��6w�㐹��k6"<s�)`��#�(�'����&�`��ʋ����ø����e��o,���؀9N�ڵ�_'$ c!��w=��˹,��ti���I`�g0�K�	�/x n���B�Up��'�\���a���1�Z.��:<l�W��J�r��2��.3��� ��b���W�ڍ��!'*6!qruNO�aH@p���D�+�R��8�A��!�w���v~7[���҆�q/3�z���ь]r��O�D(��Gy+�'ą�o~�4p�t�3L�U���B/�R?u��2��g��q���(^7cD��#;?�_`_�&��'ޅ��{��m���&C��C#A ��'1����]e<���&�[{�h�"I��.:9r���ۄ'� >�I�8�E@nk��)��C�r��D�p/��+�c�ȷ������zϮ��.��u�3�PY�$iې���%�?Qz�6W�pH!.2Jc=Z���ݕˬC�jHvg�r!=J@ы�墕�>������F�m�qW�Y�͎�bO���B���5��j9�X�.��lQ	9,ܪ�Q�Q�!⃶�4��y�a��.��g{�V�'�1����D��2�H�ˤ��=�\3x�J���u���n �����Hn�LP��f�-��Z"�m���C��2)Ϫ�lp����EZE�I]�qdT7E�����B��l� ����m�p<m�!2.|��j��-�ښ���4ʹ7o�-���L�*:�	k+8���zxSV�}k��4�nn�DYYYoh,�H��"��n9�hH���<��q�p�q�"�w|���I� �	7Sn���G43�蝤Fu����k���/�C��p��~bz��{��Yp?+YW��R�ދ	�%���1b��(���62,�ۅKq#�C�(����fO��_���\��>M�U��ͨ���}>�E�߯_����Lh��NZ�~7{�h(�V�������l{�Q�+C��Q��p)S�|��_M���man���&@����R�՟���Æ7����V��tgTD݁�^OG�>��0�0k�H���2�&c�_CgL:"x��p�^:�f�v~(\v�Y(㎧��}�CZ�����_զ�8!g���΢��F�ۂ�A�\���~t��� �!��)-�)W6�7"v�ZH��L�A��������7�:H�,!}��c:���o��>�R1iJ����p�S��`=����a�8!��Г�@2�8�!�Op���ơ�ܜ��0�`�(m���NԮ�T,��֌H̜��~٘�l`��e��7�����t`��/��x�G���]�,a��4w��0�0CjĜA?�EL���b�w1䋞Ӓ]br]Q��l��<ζ����FGqW6�7��܆�u��������=4N���'�ǿ�Z���ŷ���K"2�)��l��_�D\�G��%��}m��Վ��7ҧ߳�P6�f2�%2�*���G<ޟȅ)�;����[�s'Y�#�9Q�W Gsa��Mjq5n�nXࠅ8��^#�Z-�� `�J0x#m�OěA�:��)q�i�a@D���=�P�Q�pj�]�R�j��A�A��"��^i���-��=�'�Y��f��D�L�N�ޡ�n�-������6g.|����>��H���L��L��&.��!�;̚ମ��2 H����tuyˑP��ɋ�E�x�@����¨|�b��/����(���5	;�&�e�G���`㖰Z�xl��&SA�%�'(�|���ĥ_�P���Rީ�ݲT_�OJ85c��\Y�t����b,���~�蕡Ϙu������Y�W2~=(���)�AcK�K�G����uݾ��b����������B�}C����	��'�C�Z�Ï9��2�\C��#�, mx���d���aI��6�r~ڲ>��.P�_�{Ko�G�GN_ů2ls0� %��x���}p��_ٕ��3��!�٩d̬G~O.&�������hb���B�Q�^��l;�05-������L��� fٻv���n2sg�v�.E"���j�=��~6�]�A����_x�v��9,I�d+&=n4��L���:,����S�i^d����*��5�v�65f�i�`\	�����a���ovXǹ@x-��Gx����h��Tp2�&�ujtq�i@/��3u6���\�����½�ᴵB�/���k�;p�Q�?u��o%쨘#���L�JzU��wQD��6�\{�f�ڕ��44*�  ��3��T��F&�pW�JJ
x��I:���}��$,~�2����s��bt�!,�w��Ѕ �{��]���{?B����N��!"�g�n#'�-3�\xj��@�`5E��k�����j�;{�?*s�t	-iݗ���dʷ����~�{B�ō�_n�T2���5%�-'�b���`�^k��7@.S5��N�}hQ�!�G8���ӷ�|3�����vsj 6�x��B!�@��L9�7�cEO<Y�tlG��O���3˷{�i8n�.>��'+$v.���c�e��*OW�1��4�,�9;L��0B%4&`��f�8t�9�Y0#�09�|��j$�J�Y�gwb�p���h��j��^_F3��G�R4�;C� ��v�����x7�FM�Ҋfmn|SZwWD{D}�z��
�
�$�^���>Z������:b�d�$-VL��*213�"�F�s*!���̒A<B� ���k�$�����t������8����PO��R�N4�By�����!D	e��0p���8������4�V쾮w/�1�n�O>ĸ�a4+q��,-�6�e ��y��%b�j�nK����4������Pc�ž���d`z��B�
h�b�2��E��,�X��[l��'�����z{��ws�:R�:/	l��0syz}a��ty��=�ؐ�6rىu�yF�+th�(��b:)�{~��D�.�幊���^�B����h��'�}`�ym��+
��I�}�8 
�&σ
w�ޫ=$T����W�*����p3(�V�҃�)2DE�0�Z���	$gR3���}&1@3.�����y�I����.gtc�T���w˹�=�Ï�Si5�wx.���#�S8��J罶8�TFoQ���y� ��dk-�"	_���3��)v��!}b3o��pk��� �����5v�Z0�����y���d����GĸV�φ}&�ɚ^�B��.Γ��i�c澷���uK���kb��J
oOf��s�r���Xf"�M}f�$pY�(�|���[A/�r�KX������r�����Ķ.>51k���*�~�rH��`Ҧ>5�&Ȳi[W�Mu� �ZCn��5[ �����&D�b�~j>!�!�w)�A��vB�m�V�����'��KXVKW�� ܼΔML���[�_��4>Cې˂QJ(���-����FBkA����7%M���4B���	�6�>֟���ř� �`Ab�p^���0�i�S딡�2��GSK�C�%63>p���t��ZU���٥;wO"�������ϥ� -��(��	q�L���VD���?���������kr����nt��	M�� �%�Z��uj�|1�v��7���;�����6�2( ��0�ldv㥧��Q�$O>��/a��A�,`^�6h��}Ob����*\�bg^��>y�	M��]n�`��"ߣ+��	=�LQ!�e-?�E��Q��k������
Iw��#S���C�RyF30�q� �V��n�rDH>�Y��jCxo��v\�q��]��*��?a��U�Ȁ���Ϗ��D��F]�S�Ӗ�t�����Mr�N?)�횉_,�����Q���;:��r8����P]�Ź�w3���aj�
�� �l�Ivx���0-��MZg�޾N�]�a�k���0 0@�+��J��l��'�|��!���|�/ʏ��Ţ�t^��u^қ^�K�@[f�"�\��褒r��O���\*���{Ӂ��W����*�bDC�p�����mٙ(�3lͽl�6d�=j6L;<d�z�W-2X*��Cp"��W:ݞ6wC�ެW,�9��,�{����7���� ��M�F����I������S'�"CYR�iR�ɖa�P��2������^ ^�زr�����F<;}����$A,Zx8�=4�C�x-.�n��"��uy˅	�L���2�`B����`�u��م~�Qw$;*(���
>���.�H>i��:	'm\�[�L5t�O�9$���+e/�[\�pR�>;�V�4d�8峱�1��c�?[kl���W�9�7�(5��ޱ�X��~g\@i.(Q>��)�����0.x��V�1�3~���_C���DݩsU1�����J�1iJ�4-˛�="b��wz�w�#z����'�ѩ���0��h�P��ݲ&�ߘ�>z�v��FRU5[z'���w.�{o��Ĉ��옢�ot������|FTC%���G���QUWV���Ւ��	�>���K��[ч���������6��[������ZWa�r~G��l��Qc-����ذ���h����P��;<~��p���^ຂ뻅Jq���!�&�&�(�m���N��ӯ�7��H3��ڛ��Oh,*^�e�m>���#����X=72�zͪ��8��� t݇�d���+�0��,��>�6Pqyp��ˤ(F`I#6� �>nҌ�_M��,�Qܳfy�tv�E��âPC�Ǿj�o��f+�y*+`ڣ���s���Bf��v���	�;�R&��y�+�v�4�W�����趴ε����g�I�����Pӆ_��Э�� �uJ��2�Ɗ?���^#��z`ח*1�a�:0���S�*bj|� x������K�j�t��E�Z�'�xi��F�� ��Hvc."�u\�қ����Nx���YV��Q�0��͹��	�Y5�v0�����<DGBԪ�x��Լ@�KQ�87X�#1�*Ɗ[���3U�E6�^()Au��o� T�6�L|W��[!�H�	���� l�z`�c�ST�oW��-�I�PS���)����p�/4"���J>���SY�e`�� ���*��|�s�S�8*�s�m!;9����ga�cw19���Ce����R7����^�
$���&�5)���,'�ZW�=ǭ��.�^u�ze���~����� <��hj�{���/hf"J�Gx��2�&��(�M�%��u=v]n�|�_�4H���o�<��"�d��DF�d�{zŗx�ze#R�?��?i��i�C9��$�k��iO�P��*�������4�z��G�	�n,���#�>�v�����l�o���藰d�=���r1w����18��#뷊�G�s���������`�l�qz��a0��Pt��j�r��[��i�� ��#����JL�eq΁#� �������GhJI��X�+�:�4�<y,��؟�4�C�3�O��>�> �p��]t�c�������fުPQXb��B9�E���;��8t�����.�]?d���뱻^�Si��h>2��I�J>F��Y@?`�k^s��P��wY��K�!�½!h�i*j�#�p�����_��^!6�4���n{�pv�v�d*>	k7�*dO���ɳ������BhFg�9҂��0�j�/x$����8���� 㠙Y��N�0��n)/u�[���厥Z�#��2��`_8�A���fy!#�4�E�����ڕ{��C�n�1�%o�w�Ǆ�N_���P����Ì]ӯ�%R����<������v!�Vih���l���k�����~����l��}T�����M��61��DB[%\v�!˔���w˗2N�\�7D�9��A���K�4�c���y�O�����Qm��؛\�J����NՑ����wV���^�jc�p�!��u�*	������a8t�ã�^�um�r�+��!