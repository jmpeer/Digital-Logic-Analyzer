XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ݓd�� �׿�*:��p�+�3>�~�R��u*1Ŝ;�^y}��,����KHse�em>l�~�xh�s�TB���!�`�`�)%ߌ�t7HVv�W"�J�0��-���U�1}���������Y��P�;�&֨�ӭor��z~I���~��I�xl�?�=:�Ѫ[�8_qFZ�sb�o�%�_�o�'~(_Kqhi�������
U�oJ�*H�&c9�-��G���\�S�;NP�Ȫ���u����G�:H�v�y	��c%�����h�w�p�\����U�j.k�:�)W��(.1�Sc��{d�K��7���pƾ��s�<}�(nQ���r��"�M����0L��)@��e�![���\E���nÞ+�a��?fvW��O��y��(Q�����u�5K�k��Eޝ9���!�7΂�ru�[vʦ��T&��?� �d%j:�rd�����qm[,McA�G��8ou�R4�Nཆ�֛�Ԡ�4ta���Γ��6@����v+�!�T	9�i���'���,v��'K�H2L�N�A� �6*���	_��Sy�ݘE��j����ˆ���ӌ9��w��G��dV�q^�ɭѽ�vK�T@ǃ��pL��{=�&Z+�1�_�ur�2O�jϑ�l}h4L�w*�_������i���ꏫؔD���s���SR�C�IڋY#�Tx^�4&!k/_���fKV�(�Q�SN�~rS����Ꚛ�ɓZ�Qߧ�N(mj*�9:��3XlxVHYEB    3042     c80�.c����H�E=�;,���*�M1�`�
�<�/����l���tǪ1��D�o����V|��L�L5��t�Y ݷ�bE��wpA�P�VK��]�F�����\vx�"��6��-��is�����+ҥ����~zrt��Vukj�T���ҋt/'�����]9��| V;*_ن#Wx���z�&��Y��$)�5�γ@�z�8��~�0�\~��"p��"�|�?�Yb�-'5h��x_�p	EǸ��GOŤ��C����1Xs��#���t��p�� ���5~�U(l�0�\Z����ؖnQL�zL��^���/C��U��fQ��(X�%���=ȯߘ�D��#�:8�<�d�m��M�A���2�ފ���MU�����iTn���G=-^�-�Ɯ.����B�թ�IY��M�r�Q���r�<kg��V�7�b}X+!vj[�e�� �����kl6`����FA8GY��mJ5兵�#x�٦��n"��r��	Ϸ��}�ԧ�.�һa��Y�|��>�N&�C9(��9�w(c�-?���a&�?���gT�x���� 5Z��:ܻ��JAm{�P�03����||���u~>�!�4��q�����տʺo�7�`;Y�_����.�,d�T7,�h�/RX��Ӱɀ�w�f�}1 g-��֔���sl��"�y��Ϛ��z)���u*��C��A�nw �q(tN�Tn���i9�u��/t�f�\B��dR���1��E��ho������s��Vl߇e��f���+J����j�w� _	^������1���shJ�6��(�^n��K�|g�i�,ư��̣l�6�W�8�n��8����x(�6S��9P�&}���j���^9�e#�qP����*�S���"��/����WFf��޷���0�2p�@��=��s�A���R3��<s�&wv굽���^��#�[��[�ێ��v�۴s���|�le�@g%KO�m;��2��dd#H1kF�h�#Q�y0����i�}D ^�A0o;N����^+|���e|�=�r����h���<k�|���^������;� 3m�Dm{�$�5;��aU�y0J�٨p�c�9�!�g-��Yh��#��X{�+ � �W�q�X��j��t���ա]!�ê�MG�%���0�g����c�}/6�JZq����t ��� ��������/�;�� E�F-r����l�hX��k��C����#u#&{A X�e:
q��.����?����6��4�(2���ۅq9>����%ڥdE\aC/���? ��}�c�P�S4�v'[,��"����o�u\G@&��fA�|GFɨ�c�����#)�}.��[��u�snjYQ�����ˇ�Ov�,�%�G��b�ro%�f��ˀ���C�A��p/�`�(���͗�c�CHs�8��f�B����!Yt��
u�������l�����^_\Ƿ���L��ۛ6�kG�J�A���+t�>�����|����Af����t�rKz���HP�t^K<2/��}�؝���r*iƟb5E�T�.�I�Y,�>iQ�HM<YE#�03�����ˈ1/�<��"L!䕉 K9"�R��5�'W_�6��d�3kF��\A�X��{��{�t�g.4�a�i�c�劎j���\���6P�";@����� \ro���?�P{(��cn�,��2�=Ƭ{sM�a���OXL�{-|B��,IT %5`޿T��,��,_P�!o=�Z=��ώ+� �m6H(̓b����+bU�{X���
��S��ޱh*��tّ�T�H��:���,ku�$����G	��$� ��)'�yY�� s0�	-|Ӣ�8Vs
�<�c�Hd,���lש;Aq^�׋�� (H���b�3v�Nr/���wuPTN�$�y��5�hc���ۧїKZ�f�����ɰP�A�$S���c� ��I,�����wB��DHƬ7�,��7�c]q�e7�a뾀��J\6t�5�]�~��W똹�{��\�������+��"����΋�!(ZC�����L{'W��A�NO^��8�*,�؃��X��Π|A�w�%G�-��`����)CVU����FՈy{W	v���?�ɐp.�n�Y�(�����ڟ�YYVJ��&%Aᔣ7	���ߩ�xo�u��X�ʱ�� ^l�����=��Fs�����S�{��#�-AK�4����+�	XQͺ����e0_rv�[@0=u�x��EJ�p�ko��s��?��U%�x?x�Q�\i���Ű�\�g%tjw��9{�B���V�W���g��!��D�G�S��]�6�(��$d�DD���q4��]e���E��L��A�r�<�� ��8P����׈��Z� ��m0��;m�'t��J�iO��U���8���PM���`��G���
�Y
�������/+����U�������4'*d�_����c��K�'�_��8�S�xj�����E��*�2<��/Z{�N���=�YǪ��)`�F����);6hH��zF, �Ɯ�P�~���W�9��A�����(p`�꯮��sݲٝ�-B�=���[��#����W.1�G�g+�����,�=cz�z�lh�U�`LZTz��C��)�c��Ҕ#�yD�����px��S-M��n].����3��t��2��*3.E�	K2�{$ |הA,��U�\��M���)��A��o��I1dc��/<�6��/�/�c}���߹]�)�l��b�H��H��H"�~B�SH�� �r��tP[�@���r�:ͯ���g�dyu|��ۗK>~��o}������de�rL��_����N-D9�fK�0o�9���μ?wE�A�tǰ�����{a��5�tMbW*�c�~�j[�X$6�5q�+4�2u_�9Ϙ-�U9a,4M�!)�)|oܿՙ��Sb��s*�nPi2�JɠB�u��N�mu�E���,������i����H�(,���C��(�ΤQ}{.*W0��j`�O��v�k��]��23�.��G��>v��_q��O��14���Jn�YM��g�G�)�o	�b�k�	����a�/3;�Vv>£ā*h����}ϣ���u�k���|�rL��Ɣ޽4U��