XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����n���X����l p��W8�/�Dr�������5Ñ�N7A{�g<����,%�'N�j�
F��2jܰj���QT(#�|������s#��/�:��r��羹�z�Ȗ35)X9bUK>�����3%!������fp>�.J�&�MbdS2��X�X?�IA�"�����Yl�eNEL�yY��Q%��?ͨ���X�"$��d����C{�U�^�s&��_lv]�S	�K!$P~�ǃMxCgx:ޫ-a���GvK	)ۋB����B�niǋd�j4z|8�>�Q��o1LD�>��s���#�wJԮ.�Q����{���`��}Σ�ؗ-�U��}�罼Q���v(5�an��6y��N3���t��.���[�$p'�����ٿ�����k�)��P塅�/��la�\��(��E~&ͅ6�"��/��gS��(%h��Fk �9qg{R�!&!z�����"oN$E��{jܧe���:��L�U� (Vf��$~��2T/Z��^�@i&d�!y��Ț�m��P7�a��4�*b�JO�lR��pFe��P.�� ����D�%A�H��c{M����SҔx���e%#6�C@l�桙V�sJ��ܷ�h��<Ok�7�)�u1���('f6���@v�zԑf��Yv6ڬu��<'��Q��9(&��Tz�����D�K�j@���VWMp�C.������Y
���m��0�ё� {�h�����2*��m�^�)4L;ܯi}Ey�'9xrCA#�XlxVHYEB    9732    14d0!��)�H2[�`l�!�[�Q.� �Cp�1sHbd��X�7���'�O<�
��Hg�K̝q��[u��w�Am����C�,_�:uT�lm��Y�bڜ�1��rJc����B���X^^ 
�K�r�x)��NZ���e���Ƥ%��S�V��Ҭޭ~�(i��������<Xq�}��XL�_T\�`�6�k�~��`ӽ���I�����q0�i��|� 6Q���Um7�Fuv08dR3_���N��^m#���&=M6,�-<��iRk���!6����	Em��H�!���g���`u{ޥN�!����?J�z�a�w��D�l�����C��=N��u�y&f�Թ�����z���<ˀ=�W�	� i׀pF^��o���tڱ�uawV���(2�����2��T���W�����vŜ�n#�fz��Q�>z�?:�v�/$!Tc�b��S]G4r�ԛ�x�g����?�:�cU������#�s���hĿZU=��-�j	-��l��|��)ɪ�[�qb�?C�	,�|������V"DC w�}�A���:4��.�H�9����h5��Ec�y9�C�p-Ơ�9��˨A��|�"Hy�?�ߪ��z�٠�o@��,[�C�p�^L�@[D�?p�v_�|��c2O�&�{<�% ӵv�$�)�K3/���/�	G�>�,��zB��>v�^��`��PR��Ñ�� ���;�F�V�]���BD I�{�	J�)0�)�х螖e�:�RW>h8*j������Uk��urmf���%�*����, �N'%���f��~����t��<0��Za)�v�M�i�`f+QiY'�̸�9N��I�t�9h/]sKg��d�S�I���װF �P�2�*��j�.eM����R[����x'au�M<�~x�u��;	Q�|f��$�B0�_�)8�����d��O�_ܶSrТ�y�m�GE��Z��:eSqԜ����b�	C�|<Zz�W0�)=1墋o���9c�*�Ca���l�����ǯOGh�ڼ�z���M-qd��̉f��߼�]ޠ��@:������TR&-CE)�}V˚��c�Lvn�[P���`w?�f�q�C͛}a����ճ>��]�����5�V�cI>7>q!�tپ���b�t�bHmD;3y aL�����9�[�[26'O����}�B��϶�7�e<T��\�b9bIȲDս a�١�&���������v����`ROO��t����+ݿ�Ѩu��0����K�a[���^]s�N�nt�bK=��Z��,t0L�@��}'�� 4�]�z�~��~��~=���"��OC�O��02(5	��Ex*��J;41CD�X�s��'�*PIz��/r�p�:�XV*qB��Igu�!�X|Hc1�k ���v7��>��->�KrQD�E)�pᏍwx�F�p}P�윊y\��
>F�6�Ъ����?lyB5to�=782z� �f�8.���DA	 �<�eש�ʻ5�yc�5� �ɵ7��Ss�.)���d�w���^2�j�-�+��
�wK#���CՌ�<�����j⌹��a=��/frn�S�Ixgq�<w8��3	f|��X��N��AB�hr����s|p�k|V<�HX�	�ۺ��]�ѭ�� �#tQ��|�F�s�C.�e2խ�yP��냫��h]tD?� �z�g���^_�oI�q5��l��������!i��&�o9�5��O��*��nE[�W�8B��t�}���\� �"낚�6�%��X*���KQ�|fK�P�P���FP9H��c�jh�mn�p��{�j&�c�Cݕ�����@�m��q��Z�0�Mq{5p�yr8��e~gף��澂@*�
6j�<)�5�@��Kݫ�v��Y�2��"�.�6S��?G���3���u�֊���� ,�|�fL�ɩW�V˗XS�A)�11ymK�b|�!+e��`�T�B�1SG�M>e�4�_���~�'	i*�Yó\U/Й�ǉ&W��[�
?� Rf�}� �X�V&�������`~���h��j����On��0�]�=?���!�����	�M򁽢��5<���S� ���.�Nv�7!{�Ѥ(կ����'��#�wjh|8���΂��2�6��7>Ƴ�U���40��b��`W�����\��<�}�6T����������]|�2�2����*�5��?Lt`�Z/�8f�ƌD*�@v��Z�vy�,��/�?�\�n.�a�_D0���% Ch�Et��h�,�*����C�S��֕��h�d�6�@r������8�(�S�!�G�kl�����b.+��h8��R�lH��h��Z������,I0�cv��pM*��d=�x=�2��$����Y����1YTf�z]m���^�������4�l��DnR�"uz@3�����'ܵ��J��K;�Q}�ɘ��8�5aS"ݐ 7.$�3~�(e�Wg�X)/꾧,J�ROz�Ʊ��X�^�ap�R�v�����-�K==�E��khg��f�y*�b����=>>sJ��j��v}}���&2H=�W����J/9"u��ys������.Pja�DO�q� ��WVG-UCK����3����@]'`Ͳd@WT��T�����O�2�_�'�Fg/KwU���(�����{����jz����F�
�@2���M\;i�>w�B�=��2�H��s�c��l?����9�i�F���%�6+WFy��G5�eu�x�������*��A��L�@�1����Iz��j��9[���o8F�،F�L6�>���}�O�ᜌ?|/l�y?<Kswqm����'����C@%C�\�;(�b�X�f�t�혧�R]Gܧ[44??�N�x�+@�t���V{� a�%����G7�kYq{f|�tݾ��Ħt���풲���n/3���iSۣց%+���谵�wv��,�L��7N�"'8��S.R�2ة��q�D���Ee��X�v#�CeF��@��9��b,�� \,6F5~"ێq�E���"�+�U�`' 7�R<ܱO���.��b�0���BZV8�Q���4�ʋ~�@/+����Y�u�pU�����|��a4a�`B�qx�b]��#9|(�Cn�|t�ם��e���V�xƴ��Jԛ��ӪT��&Fk���l�>��z�G�h��)${rK�hl6�W��c�V���Hiʃ�0����z�7ե©_13�=�̵J�����|wZ��H���W�����O!>V�3'�?�#�M�"p����ta�T���vn��p��vuI}�>���=n��%I6�m%��e�y���2��ҳx�'ݦ�^|�<x6VX�q�cC|":),A�?ϝ���%/�靭�6T'�G�ż�{S�]+I�h8��զ��iۣd�VnC�uv�[�~��36�5�<��$�t�2��b�d�7�H)�>��E��
y��QXkVX+��Av�;c�wyޚ\ABP�����l7�����I<��Z4��ܺ}���ݮ�t}v�� �A|����O?X�&��g��cf�e��������k#����m���N��x�K'/�^g̔.�'=�5c�x��<Z{w5^[�*�������}����U�2k*�����P�u���>P��S	�H٩���}c3 ��lj� ���P��sz�ذ�Ba�>�^��8�_��adG#HFG�紈A�;�LT4w�
���l��B(y����r�M��g>&�%�5lm��\��L:.u}�p�9{��C����/z7��@ʥ��9���I`S��L���&ᒦkk�S�T����?`@�QI�j]n�Jv6,t	�'}�������U�C�Ic�*��|�&Z��S�<F,�֪�\�Gl�i�I�� {=��x�|X')�M�說�6ݏx@�W��<unt
�%�K��
vb��T]B��q!h�E�X^����v�AJ�P�������|%3�~k��Q�c6l5�C�jpK왒��$m^��C�*�>x&䇢Ư�u"�]Pít|�A��xE�q���_��3q�]��N��D�;`\ �fbw�3��^�*F�iw�۰y7?i0R��#s�npSF-T�u���Oq� l۸�����p���~�܆e��}�N"0yFO"o\%�O?�쏔")zV.���RC�>U��9����K0.�@Ǜ�Bi�����R�����&�,:���%������sO�D��e�A*��ߣ�g��;�9�_"Ez�D��ve\0�f��?�;Bc a��H��e���VD�WV�,�B�C?�d��|w����N�Q���@!X�t{��h��6��{�wY`�Τ��.���*m.k;�`��lT�W_dr���f��<v>��Q9�w�N����E ��Ũ��f9�^�z��G�M1/���=$�/'�Xj(3m���=���|m�T|�,��\"󳘥',�]¸�\읉a8���v�k�1�h(@/�rT�4y�^R��K�f8����}�MC'��c�6���M����c�N:��mFX3�A�֒K�� ��zk��b@�����"�B�)�� ��:�����PJ���=��:�"�B��-�n	��f��!%�m:<R�҆�F��	P^�HP9�hf��Ұ[3܈!�X�H����bޚ��L@3�������I� )'�jY?y�x6�!�\���eS���H������V�S&����;�R/(%R�;7�2���G^�*g�"�F����b�t1ƈ/���Ġ\�w-�ڵ7���o��sDӪn[�w�V�T9(ET���2_1y[�`/X};�_!4���9�j�Ug��,��^����u>��)���������.��%�v|��w���S��p�&$�\�&��_��&rÑ���6��YxS���&�ba7�����\c��p��������KM[��m���;B����-+���� #���'��9�%e;��3��X�t�xI��_Q*�6dk���������Ft	�--��dȓ_����P�*Ĺc�.�K?��8Q����(�O�o�rL�9g[���(v���!�)�^����v\�ax��}��>YV��`�^l��#^�R`����K�,#f�Hl��GD��Jb�'%�k`G7>��g Ϋi��U)!� |Q�M�k�.o�h��	��;q��,y-R&!�k=��s�T���p���(
�y���w.���Fz�����Z�b[j���ן�+����D�tQy1|s�߂�0Q͈H