XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���x����v���Τ���ftŘ���������Sw�[ �
��K��8���+~���{��Ի���6�]��]����ㄟ��xW��Q�+	��<r�64�� �dE=�k����rK��2���N۝��dCo��mC�G�v���2e&�;Z+C[ϙ��1��Kz���l�R�U�O���"���/�6��ES�2,Ɲ{B�C�w��k����\OB��1�Қ�7Lk=U�g�)+{bB����fM�7����&�����`,�oZM��锎0���kk�,�M��7�t�	l�S�UF�vx���V�F��։��y��<�2s��} �����YA�?c^o0hL�D�B|��~�Ƶ}$/�|�q$E"�^ҿ����e�A�݀�HvN��!�Do��7wv�� �Le5�%�l��e7h������;d�|71
���

Y�e�Jn�\�3	���&8�`����0���xl�/j�wt�	��z����|6�����]�$�B*k�E��;��5A�13��sy��[|=�^�.8ݛ�̕P����G�L��S�ٜ���NO@=�Bi�B#s���&$�x�37�χ"l��C("�j6U������R�l�>���oÛ�U
Q`.BT� =h~r�fA��C	@qB��D_��e@�"QP�Ƃ�ڶx�ȷ�CT�S�=;���=��'j&���PѬ�E8�D|�b�P���U�5Ms��)�,��=�e$+]&�$2�)�7�XlxVHYEB    3504     cb0��s"
�w��	رh�g���V�s��FA=��V�7T��o��]S�@C��k��=ʂLq_��O#RY�q���US������Z���o�ͣ���%�²�}Q�f|j6%6w!�w�e9�y?�l-��E^QȬ�!�|I�!L�٣��:S�p�Is7o��q����b��Y(�Cٴ�|�6\%�ۼ�I���.�K&{�eK��v�_�G�7_v�C��/M7��ƴ���Ѽ��ۮ�A%�����:��e������J1+������˞�8�d��y<�9&�7l��<�S=�����m�Զ����s�8o����Ļ���e��`.���2βf`HR�g?sZ�Y���++�Gue(���}@\e�%�y�p�d��h��y��I��EF7Ƌ�1�	�tN�BuUTi�S�x��} ���{�-Dq����U��o����9)���3����>9�a�GR����;;��f�����Њ��j�9��= �e։#�1-���!N�����e̚��o;�Qh�k�Xަ!΢6�<O��IxH홊���@X9$��f�`k��&k�6<t1
׸q�u�n)�	�t4Z�<�?~�f(�P��ǈ��;e^��~6ϓo�j!� �^f�F����2.ꉉ\����OA��(BW�y@��kkU�ٛ���TΉh>�P�w��`[�x�ҁl/�ɒk���I�C@JH�������5N�؆{а�7�ؙ�x<�<N�O�T�U��G_���q�gS;}N�%�"|�r�Ҕ��APJYAOkm����Ӑ%��� �g;��{����x��]$�-J�L7I=w�\=|�<,�8.[�y�'C�)����Y�z���_,711��=�3�9;�W���eK:�hq��w��動P���N��n7��J,p�
��Qt�N�o�%��a�:�o`�`�q�°��[(Q��L��Os<3	�F"��p�&���g{�D�LЎ�R]#�1R�C䴜��
R)�����t��C�$�::�k.�>>��6�˯&��τI'�N�/P�9z�I��#��i]- ��@,g�{QoXY7�� ���;K_���|5;��ͤ���j�V���r��sʛ�1)��!���*bE�@�o^淩����4�>F�`ⲗX@vW��Y�&�BC�uF�����@��Eb���Z6��k��n�_PD���\K��Ǧ��F��b��8�G��Ҳo���$>�"�Ì���nN)��f���������Y�(�8H=��RLF$�Q��I�q�f�i-�ܭ>�tf�4���jabV���WlǑ�h���r����`Ɩ��e&0� ��n\�;��o�y�9���U��`���V6p�܃�K�BF�+�r27v_�;��qØ;��<����n]W�f�t��Һ�?v���ge�K��j2M�	ð�HU�Ԑ[�> A\`���:�m��X@���Bh����\%07^��5㩯5�'RM%^�-���k�݉��y���:�&�������3e[km
�K�j�M#�;�l�fh���VVǆKg�{z(���)F��L��d��� Ŏ	4�O�F1�-a�n�"��H�ʗ�y�����d����M�K�$xc�x����(�֖);�N�]a��e7;�0�8
!UR�����ύ����^�a���ļ�~td@P;����/��<�u��`�j��Ǹî�I�����2IJ9����ҳ����;~7y��#�5G�s�!\Y���SK��Ŏ�z��`[84�ܪ��B�ظ�;ǶB��=>u*�o�k��Ԕ܈:�i�3Is���v�a���٢j��.l�o6��kր⼯T�a�3����g��|���g��{iɆ�y �B�QQQ)���F��5��8JSZ�U���o5V��'�K��b 9���M�2�<����~i*;M�[�L(�*(:��'n�4̪���.�2�����Y�&F�&<�&��3��b���Υ��������t4�S�[E�oV�:g[Ύ3wi�c�����ӥ�	���@eʵ�	��z�D 0�� �
�/����6Ιq��&��B4�� �$��T�]'�p3�&X{����kL�ʫl=�3����F��+�
;���#��
�K�v�Z��U������ՃA7��|Їo�ҀSe��2�޿���d����`k�gw�n	;h���_�(�36����/�o0�$�K��>V� ��y;5$БM�{O�2̦p2��/3��$���7�����ɯZI�<[��}Bq�Z�s;�Q��a�e��M�Urg�����oOd���A�� 2s J����y���*N%a��x�LP�d�Ά�#T��Z+�6ֺ���2t��!�P���h�� TMjY�D��{1�qX!� Z�k8*,��Q���_����J�L���ߓ��
�J�6oR ��/\":G�ETx�c"�G�ЎV�Q���ynI���=q�MU���1NwZ�d��-7E���x:���}pmW�t�sC�f������.�/�-HX�
��rc�����< ��w���Z @Z	�קXD������,ke�ə�	4�]~ĥ�C���=��v���Ky��4t�ZbT�BV��A0�=�*�e��;xV��2�Z4�N$3����MY�r���J�ߗ�5R��RUq�i0�'�گ� 8��^F�/yxrۯlW2����,l��H�$>����H����Z^�l� �ɖ����}.�9Z�V��UI�@;��0�M�2�4��{�Ig�_��أ�BM|l[�Y֬j���H�x��|��%$�^7���φφ�n��xp���)�Xy���hwT���4��6QL>���6�v��'gB�4�IQ b��d�ϙː������1\���sĹf�`�o��E�-�֍�jhτ�X��Tp�9Ov�T�vsL��i��gwřNx+\��Z�o���)����5yُ6K��x�R.:�PaK�����n�<�'����%�J�{����
oC��x��Ѓ\�&��1 /L����D����i:owQS676��+l'N�a�Nvr4�	2Y�>�A���4@)�
�B�R� �%.��f%��3�k��k��q>���o!��EuC+)o��8.Se����J��=R��м�)�/Px�ev85���Ӻ�� ы-`+ ?V+V�  �
��0���e৅Q�^�#y�9C�:k�YH:���A䷯�S&�t���X@�0�g�.b��%ʽT�