XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���[T��4n94\y�u���YjhL`�����HѺ���L+�yݬY���F'�o'1�l&��� ���<ٹnm��;D.<M����%�@�B-�q1f,���tc�e�h҈-y�-�C{�f��R0L~Ar�]��X?��<��1l���n��L!f��GO���:�c�~�@3�I�p�z�L�N	4mN� L0�&�Ϗ�=��yְ�<�{I�ۊlᛁX:����)��c���l�Z ���Z�Hg���h_̷
���,�q�4gP!�����(�E�1��T.�V��2$�{K�
�0���b|��x/Hu��F\�N�y$�ɟnxC����/�y6DO�>u�w\@�sn���V�=?n�s~2���i9eB�b���o��@90�ǨS��_�D�Ĳ�������eC��^6�3HD:�sh����g	̑�J��챇�jF��8ۺ;�;�19h밟�9����M5D>�/ �/B��8�3��a3�-h�0C�Vh]���JMGE�i��F[�Q�%���;y��Apѯy�i��6����`�e
yP�݀w���"�*jQ�S����/ �<����Qw��v�*o��$��R���K�4����a΍7�r~�o߀��o�� 48�
j���U�?�w����ۢ��s�Qjw�A�/�֦�x��{��&��{h6~�<ZI��a����|O{E���{�ixXg���bڃ=�Va�d��=�5Jdx:}'��ܹN���SI��{^�E��bq2��ؚ���;���R�U��s�:['��XlxVHYEB    fa00    2d60]5.� ��w�u+�!X,jD�r'���c�0 ���L-E�t�4������2Z���~�ǌ��e2ܜo\WF%Uf��H�z%A}��������x�-�o���h~�x�<�ŕ0-e��XE"{qR�*3�:�b)�'�Ʉ���z�$%R��T
vX�fp*�o}Uu�
z��y�9�`pT?���eQ���1�o��D!�(��I\�n(L�k7Y�W�?-Mwt�uO�J�2m�&�8�r��Rv�ɂ]��"1��~gm�� y����5n��-�&�������Ƅ/P��qN>\��n�*t��a�9I��ż� _������3���0�/N�̠���u�g�����P](���J�;��zR�W AlK|�mV�x~�P�!�x(�^����~�T�����i$P�$Aۙve�&�%�%x�I` �.�,�y�qʏ��2�X��MMX��MD��W���x�@���&������M�����
&��q)@�����s�Tf-ۃ���խ�Sy}9^�_lW3�0K�NW�)�3��X*��'P��qu�b�ҹR�\�JP��e����o���mҴ���QH0�P�r�:j�t_,�U��^e�8� ���LI?�c\��Yo����}{����b��ݱ��h69r�f�+՗�D55F������ �3^�p��fyM��@��Aj�y8�wT��k�O��>�ڟC����<J�Y`�Z���`d~�1w��ĸOM��G��i}����Q/��c>x��Ś�h��e�����x�6ò���`�P��v%����̴�(6a�(�mZ����z˭vT�yp��E_��^��J@<�#΀�[c��M9M���!݇f�	��ͬ���Y�sQ(ݿ�aܹu�M�CrP|��g.�'���^�0�8�t�b����D�|S���a���6�?��(����:�=����~O��Q�%Ço���p)>��zN��ǧᎲ`��c��]k?�V �l0Cl7�*Q�DK=��{�
����t�v���4�;[R��o����xi�T�J��#�g��V?G���>��fÌ��s��(E��ӹ���ëȗ��}�J1�"�Z�A<��U0�
,TL4���J_�B�E�u�-�2�˱��qDI`�L�Au�?jy���H\�ln���j8�#P�n�)��} �����e�7Ԟ��X�w�`�~S#�O�M`�SD������[F�����_�Y�۱.�HF
2Q
��ZE��V�����;��mT_���Q1Q-N,j�Ѯ3T��Ba]h��Z��:�3)�8�}�k�%������ing�.��v����|��)c��}!\N^Y�;���6&,cʉMό�)獰a��_��9�l�*��D�ax_�Q���S�8 ? �,�i3�G�-7�c4����5�г1�n4^�႗!�7IS�ߖ��E	M��Y� Ƭ{����]�Ć�ʧ����U��?NT����J�m�)���|@�~U��%�Wp}mA�����Buo3���W��s�/n�1�;�N�-�����X�5?Y��{��\9�e9�J��h\�:���B�,,�[C�E�_4^���_5��f`b�pӮ���#���}�0���Y��i�<0��De�3q_t�X.#�'��ߏ�6|�_����2�ׁ���_�A�Yy�O�>{[��9iR��9���5XvǦ�΁y�n�xN�x�(�����i:.���Y�����!�-���ۏ�#�uT�Œ�&_-�된�zϪ�4�_�5(�����`j_���I�+��'�
2J��҃��k&P�r����*�"��Y�Sqc�	Z.4;��&%f1Ҡ%A0�m1)����f *0o�7���%���Um�ţ��g��1.�N��6�r�D�&��9��3���nGa;�z+WJ����l��Q���?y�)ce�u�'j��#K�m��f��.����>=!�+G�Tm��ݵ�!�5F;b-��_���f�����Ϳ;������ǼU�a;#�
�ꄏF��C�#��n�P��N������˝43l��1�������kj�-IDIU*D(�����7�m)�}LnZ����n�jHp�N��,�|�7~,��5�W��U�wH:�#hDF�K4<~�gM�����	qV�xi�^8S{Hˬ�j�L�l��C�)f��i�Ep�9����������#��	���Q{��=Q�z�4opT�'�逜�|�qB��7/�@��A+. �^^�����z�>��\��pY�>�m�:��@�a��8��Ca��ѽ5���7]?���/�==���m����V�%�Ģ�c4���B��v�V2���#V<+u1 	:<m<)k����\M��)M,TD��J$W#�� �v&��b�b;M7�fl��m�{�~߻�P)�B.�E��y��Y杍m��v����`{	�X���i??�#���ø�X�E%K+��u�[�5��~�������t���X���������鶃PTF�L¨�����+���t�0�1���',�+�@�3Z��/8��q^&	��t���S�7��i����.�o7�3ۯ�e��F'fku��q�6^��S�Ӈ[�k�]���Cqsjmh���ꧡP&���W���p��w���WR-o�'�R7eg�m��ִ��J����/����XN5��){e���B2Lb�|�+��3��|���c�_"S_��G  Ƣ߭Sp�o�,GY��('�B�a�)��< �bS�8�I
��q�{���o�d������8S��X.��Ru���r~�+��ڰ��x�=�Tf��lp�v��k���s]�EXPYZ:7��(������FDi?8p���9:@�|��������?��=����^�Jb�]��H`W��ۙӇ�"���H">�	�2\v�Kɕ1�!�":
DA���7eiU=E3F �K�X�dB�{�6��v*��gg����S?��ޑ�]xҏ�8�(���z�=�\8%��B<�����,`�v�j�T�n��u�	������d'��|gx��ȍRK�S�����1a��]$�ɃJ�UMr$���Hօ$�(��i�H�R���;�W �&�3%�.v"w	o�:9�"!0�E�f����8��̴��X����-:G\�k�r�]�=�Θ�6�-4��	�7z�Ϋ6X�(GPh����/�� u���ك�����:���� ��jO�p5(*&���6�{v��i���7u���������k��bsg�@6�:&�ɪ�T�i��mSnT���(<�����?����3�=��Ȩ�V�P1z�Kå�/��������Q�<�yMg��%������X_l��%��x����lŁ��t��f��d����{O*�k|���%�id���~��TB����
V���;N8�'�7��E��Ԅ��e�Aٲ���׊�Փ,F���s���Fm�0�J���_�{�fZaޕ�<���X�'���~v��"�̋�� M���[yQ��g���i��k��p�g��x�ײ�ɡ��������a?�Ҧ�e�a|�H���kv�wmEgSjz�aMW�C:�ϖ?E��#�`�wh�q�$��ԓ�X�_�k<�R�ġA����^���A!�K ü�q�~1������ԜH:�� ������P�� z��f����Yr4�Y�n��1S�{�z��M>)���E�����i1�:�J���OImiX��i(&
Û$�<,ی��g9�o�;.��]Uf[3)�Tޑ���f�]k2}�Ӱ�P
���~Ŭ����;�6^_p��+_�1~fgE��BENUgP�@}��D#o��"l�����Й��V:��1JĦE�Ǿ~��ک�vFNc�����\�f��h���?���{���,���Z���]d�^��⑻??T�u���� fsULj�E"�]�� Ӊ���vљ4��m����	�-��x�KQ����[�c�ǀ�e�����7Vr��?����2H�?��@܅G��?y���S��I&�⠔��x�R�g�Sij�_JWP�|�!�K�2O)�7䅔'��t���Qo�YkLc[��`IEf)D<��Cy�������p���P�|QM�eWxPaXI�]lv����jU�qe��ޮ�:�3�>�F�`�V�J´���k�����9�`t���m*����=%8^�E��ř�͝+����,��n��� ��\�8�),��6�)��Ӻ��CB#�P����)|+9Sv�&�q�˶݋4[�+j����_�o@ޚ*�������^�9����q��FX����rFs-�JuS�:3��P�A<���>1�$�af'��٫	np'ff��%۸2��p�������#K2�tމ��,��w[��\��h�������^k���O10Ы4��_��Lp�xg��G��'yqO���y
�
9Q��A�B(W,mm��U9T>9����$��28�|��~�![��$60/��o�^�����ÆF��|����c&���Oj��s�Z�;��%1hmd�] c��au���Ws`�M]�����b�c�����c��#v����%�wN�*��}��M��ƬKɩ�<�{EC���o��}X�5>�'ҥӌ�*� �]M]�,�O[2�0��=4_�(�s�BU�_��g5�#��i��m��E8�x^L{'�ہ\�XZ��A���6��Xt']���|m	C�pk��D��޸��ژ9ҏ�q��^�w��Mq?�1��ْ*Ҫ�B�`��rn�4�C�����tM�����;90�����1��ō7J��dF��.�*K[h&T�״?N��铆���X�e:t����-��t��q_ۈK��Z�ș �DS5�Zpd���C����$�G��.���+���ڗ��Ÿ��V��T���G/{G�K�O>Oo��mg*�Rt3��:8����%0����$AO�t}۷'I�2cSp�rB� �,�lxAܷg��kb�M_� �:c��kJVæ�vgnv��Dy}�S�� ��V�q�f�ե�c)����ꆻ��9���g���y��q��]��͋Z����)Jɥ�`z�r^8�`�W$�>E���X'�p�%:�Z���F-)M�4t�36s�b������B��hb3��uy1ޚ�.�z?ư�:��#�1��%N0�������p!��^"¬{Ț+uI LG^$��2^���د�m�� ���+�θ��>C�14\���7Ц�4`.^���芙��¤���c��T�_��:�2�?^�"Gǟ��u��-x䱛��G� r2�+Ψ6Ȑ�����'��o�#~�����dh���Ti����@��i�\\g���&]2kPP��`("��i���!,�~�]z�ŀ8���z���+5N��} J���(�W��A��N�6v��9~У�.�'�B��uG��a�;�&�S�� ��K�2���Oj��O���/X���0��'ژ.9���N�ekh�q^~XkL��)��䕴���&���x�@t��g�q)�t��!A���Y�0��JX2�r�� �N^��*7���!M�2�,1��;�>��Bɹ~:�0T�3��qa-�N̊/��eq�t�2'!y�� ��Ѩ��hq�#I��>�T���n�1|� ��N�8�,aϭ����;C�D���`�K��t%�xw�S6�cG99�z��%�va�dn�xc'�$L��E���A��[�����]�m;|�EەEê���7�{���^����:�l�Z�R��u���1��S�> ӓXfepb4�Ux��*k��{z�Ev�D�FE�b�ag���q��D�X�#��,C�80��EC��)U��|���Ox�aW�(�4�22�>^��������+�f���d��`؛�6i��f�d ���d�}�T��om \#@�C��������bSN����Yh;sT�WDS�%cfܠj�ƪ��k�Ɛ.�88b��!�tZ���C>L&���z��u������!�'��R.y@���ȶ�gr9��/r�*:��S~GhIF9u	٬��:��.�ذO�=�s-�6��\�^���sv)�6.�G�z�S}�8�H޷S���o���3)ɫ0�~�5C��: �] ����������Ғ7�-��Wq_i�Cl���3��]å�qzJ��#�\琮�9lv��UŮ�N�"����),F��K4<F�G^9.3<� h����k�w/S*Q��r����"�Tk�
PG��!ŕX�O5-,�<���v��;؆;5[S҃��Jͳ��|��FO-��/�Ӑ�sﾏ/�i�b��{ȣ��u�Mk_�8ǯ�.�=����홁w,G���u�ג?`�'x�WY��P�4�|@�kϦ�T>�<[��|���:��Po�C�=�)��%�)g��%	e�C%s������M7[�n�u2}��9\��`�;.qW��F����A�OU>}�(�Y9�&3N��*�:�h|]4�7���DC\b�@LZ�728hmTHQ����ԂA<t�{}c�N֚���T��T��Z��'/Ar6������yd�P�x�I"!1
6��M�R�G&�P1�|F8���Z���h�m���&��E���6߻d������-�C�X���Xt����Fo�#ѽ�IǱ%�]�S�e� u�[	 Q���Ѫ�����`a�Ʃ30����a��<���?�mf^g¡�G.au��F��;�{� ���U��Ub^c�V�u����8!��q�E�k�o��b]V9���ڤ6/�s��{�ZL���ëF	�n��KXʥ��}��!��h�X�9�֥�wnD�K՝��SH��g�ʙS��y޶Jg�B�M�p�)	��/�O1]�aU��z�Y�dC����J��/�+�p�2�A2�sM�3���� ~$���l@r��םe���w\EV6�'3��c5|Ͻ�Z%|/���YE�j�i�����`�V�PF:�����P�_L�-�W�ϝ�-�$�؁�����e��AE싻��M4�b���Gky�D�4��cp�3�x�1��طѕ>����棨��Z�t���Iiy��2.*�G��OSg$2�՘�����L�[C�0�+�=n�fv�3��.��|+;`��C�K�.p���M��"�+g�	�Q�**ΣK�6�2?|�O����v����a�G��AZ��@C�a�����[0�V+������p,�`�,����}Xq�Պ�}��"��$���t��t�"��;��>�ó#�Qx߇�����<1��@	��
\��[�q^�P�7˱�Kct)N�b9�Ip%�e�����r�_�d^�)�N��~͘9������xk���*��N#���ݒ�xV�5���%k�2�t��S�$-&��1Ii�y����*ݎZ��Oid~6
!Vج�����5�u7��39�AՖ7���H�x-���.�7ډ�,=s0�Q 5���_��ջ��z�Q]dn>#�7'8�=b�l��q$kO�?���ǗAQk]3ZHy��Ǆ��)�xӁ�У�7�Y��ϣ.�2+%ݱ�"��}���Z'Ԋ�O9�k�P ҷ�<��\UuWf!\��9T]���[}# 2��w���M���K���#�x���T��3a�[
o�mů!�����㯒���	�	>��C����C{�ߖ��i��b�f)�Gb�C�V�Lq={��j8K�|.#A~{�N���b�`�J`u)N����&�;�$�˧J��G�E���b%w�i�-���il���I�4+�Gz��ı�a}��h�����6�vU�� �e���)Ym��м�_��:k����@i+7�N>+��?;�u���PJ�h�5��`�՘۸�9�O�*\g�<h<�CI:[�ᓊ@a-X
 Sl�[D���'B8���I8�ִPp�D�c2c[(�ݹ�݊�,w��8����Y�/�� �R ���s3Db<���c���d�:���d	�06���)5�nVwr�pK*�;3�����̞���\���:KV_<������j��8=wcq[���k䊚�yml��M]���D���<�����rQu���`��{�*�8��#���9c�+��#��R3�sj�w���{�'�a�v��B��8��Q][�=�?�Oaz�y���S>Ķ����'�S����������-Sf'��G>�7��-Ƹ���O���q�"��l�7�c�03^��5�G5�#�sb�.�fny؎Xj��'�n�b������ n�uG�tWi�2' �� c{�K7}]A���g����/��r<sV�V�Ь-���bU06�m*��v��F9�0�3�G|�i������GaM��Y�����Ğ�Zd�ES؊��3��è�yT1I��F�_7�kx�y�^LS���ɻl���ѨQt��.���lPbb�{[��{A\�����a�D
3�Ѥ�LB�"|��J
�z^m��C��@=�3���1����f6݇�N��?;�[N���0e�D����\Q�#����C���6��U�G����h��o1�nHv��^����Z����G��	8��r��zb-8�8@h�TU;@�G���D��0���\F��ڿV �:.�K)��Զ4w6l&��-���L~*.ؚ�! t d��c���>��H��I��L]��a|J�w�;���ݷ�	��`f��3٭[��"~y�!�2�T=FO����1ݻ1��x�p=�!2��2N*���W]O<�n���[�{����s�>�c�Q���yM�`���{[�#�>��� �VN�K�I����;ȏ��/C�9�Kp�͖-*|+4\ks���w4���A�~� ^44]Os��H"�/X�r���<�!��2F����W#�l,���B�z�3o�W�S���@MbFɽ��d��aCo��d�W�~�BJ¯q�0�l6	{��3��V�Ì5]V�d:��2��=�����zmEti�e��t�vo���\[����0�W�`�����8�؂	�ٯ3�g��Ekz���@�S�P@�@��6k1Ǎ�9��
�MD^�-"ʰ��» �O@�H�̤-�#��oF��i
�Yǒ4(P
��^j�����'?>+�`É�w;(y�ؿ�H\%#��1pmԺ�݄�[z:�����w��&&Xڎ�ǉq ��;�j+��ْ&�CX�D&�{�Vg�i9Aٝ3��W�13a�]l����	G~����F����ب�}{_�T<���M�'�""Wj5iA*�o+k`����tb����=A۔�R!�;��1L�C	��Q��x�x�~)����=���WJ��oFڛ�nj�������	����4���?�+@AGR����+�{H����\��tL> �i{N���9k%.�-PL]���(��̀����=�?�܇/)���pܟ���f�OW���9�H_�a�qX�`���El��ɶ!��y�C����m�j�=7�H�i������~���8wg�wC5�t.�ϓ{�dk_�sV�Pg��3Ԟ:@���z�_�UB�C�\����e���4oƘ`��1ǿH"1Vk<�=.���;)r��U3�	��"�p�[h�n��E����x!b�)t�')���q@u�h��Z%�[�CTnb�ɂ�޺�+�<8�x�Ԋ��vRZI���/��9�y�u_A���s��39L��5��
�m-���ךx\C�vY��:�V��HB'�������޼�u�2��&���Ud�f�hT��R���Xlm�̽���p?�&y�}FN� V���hl
��㪸�G���x�?|��}�k��5���Ҳ���̑Qi�M"m��"^v
�����M;��l}�X�+Ǥ�=���د�N��Gή�H
�W��|��Ky9ު|�BױH�E�%�$�[�hA����[l����8'�;�8�s���ȭC��3B��J��5���M��>%�W���	\�cAJ�,Fr�o�6�+O/j��z
&�P�����$�s�L0{�WM�P�����p,��'�`K�3��=/T�f�o��ž�8�5���m�79�{� �yoh���at�C9a�a��<�>�H<�I��7ų�T�rτ���Js�Ĭd��rQ�^T��a��?.h;c]��bR��$��8m�^�_�Ǽh�� e��V����b-&"�h�p��4q����㩧��$�����㲛_�婰e׺�o��9=[�,@�i�α���/�Ґ�O���I\��H0�^K��\�WO�h��Gq?���+���s��n��B�e�=�u�Ѱ�{P߯��ɛ��pH���K�����R,o�y���;ZQu����B�:|;J��9IjU6�1���U��HG:�oQh�E���D�sa,1@�#���-,��N� sT�ה+p1\���Z3(�[��(΄6#BUKC����S�i�l����U=>�<����R�ܱ�Y@���H� C����z���Y� w���W JZ�����ed7[^��wyr����vo��ֹ������8�}{�q�Y-��n	���6�PŒ\'�Г$8}�RC���[��Ԛa��˃ 
uXh��T�9v�e����Oz�9�(&�dcx�B*�+���pU�2#M�JZ��K)U,4Go�b�W����c�[vm���}�赥�i��ՅVP��������@�ߗZ�C���k��!�O��l�B�v����+Y[���E�e}F���)A)r��TX��^��e$���5��r�ġI�10Af�q�� ��b�����*�%�w��N����x�lm���+E��wY:�]h�Bm�d��K˺�Mv�8<��B��$!�+�]5�KVG.��<rA��#q�_�C�Jb����	��k(={�\A��+�<)iԷh-ԥ2E| �h��J��xc�DaZ�������ŗ��:���=���<��.{������N�TPSv�N^�w�&��deJ2��D���p������=@��X�P�n�E�<�n�A�[��"���p��'YCn>a�M��+�tng��������|�@�AB��/H��M�9��ЉQ���/T�NG�Y'��v�85�Ҍ��\�+��h���(7�pA�T�t0��1�i���:9�~tW�Mk��Rb���:(Y��Ua���͕��R���P���*��̘�Q��Sb����ğm�Eݾ�NZe|3��;�p^�t��23od9��yː$p�>�
c�e"F���.%��,Si,d�F5�K��wk��v��@5/�Ա^�`}�h'�b^*�����qp#r$\��]�9Ou���e�I�����6��t�Y3=ب�2`�F���`��Z&�a}XlxVHYEB    5914     f20��6?� �S�8h!W���7��lV8�_P��E>Ȧ/����^ǩ����/�P�<��EnX����?�=+/�I��j�UG�5����~;gc��s ��.�ѢL��$�ES��n�o:�;��!m� k��E�4J��l�L��S��#H�&����8 W͡z�Y|�x�oRS0�`�]�<`�5������X�s|1B�gC$��S� 3�DɦsVig$`6�QN��m����	�1��0n�FFW�a#,4D?���1k��&~x�2;���/�I�!])�w\�\�\f���=���ݥׁcd�#M����U���/H ��b[g�������w�x$��v�7W�ѣX�پD�v���3��1��7xN{0YV���M���T��/����DTA�
�>?��D��SN-r}ʗǵTԶ<�a��|��?���P�J�9(P������ew!c��Q[�7��E\~������B9cy;V��PT���=ae:!��ھ���9�Ō��q,m�l��P�H<S:7�ш9fЈp<�H�?q��G:��$j�|��A^��'V�yvН�.M�R�����F�.'GK�g���n�\O��)�������R�ATa�U&M���b/�4(���b�L�H���{����JI�Y�.�|�95"6mtҼM�-��7���<�ƃó��`6�3!�Y���\�$M��;�PA�Qc����%h�,�w�bG��@a����~����l��'��)?�
�2AI�Ál�&��`�{aVw@$�<���� �<�H϶N�*�� ��vCD�ì��1'�9�S��2��r��h3jL��em<z7vB.��&�%K�l����Ղ����tA�����;N��� �*|��?�1�ג�I��X��i�u�i���1��g���\��@p(�{Ċ�/?��P�
��<��>W�+2��g0�ת�B_���9��/��~f�7����P�gEX�Y�G�Xt��l���\�]���G��n�Nk,5�vL��`�[f" �òՋo��:�{e����@6yN��c<��h��ܡ�l�B�Z��`.�Yϣl��z5�ʻΆT&'zt��%XB��M�֍}����zqf�Du8�n�<v��<K���ݟ&Q�Ê�����C��ً���.��	����'�3U}^��\�NQz^f
��H�m��e����<p��A���H�QTe��哂�s^�z�YW��*!j����9��|�*�qt&�[�	gsYz<�F:�G|��]6Ÿ|�y�����Xk:��7��]=���VD�:�ޢGnk�������؉R����V�FC��g��=�J��"x���R@t`C)�
E[o�M�Վ�8�u�d�p�9��8�6 F����Y�ۧ�WG#��Ʀ̲���(���a%�)9��16?��q/��. 43�8���ݶ)�[��br@R]g����sO���w�q����>i�����|�O����gP��>(�;�M���k�̶��s6K��M���]S�?'�]f�x��Y2r�y�	��l�l����ծ/�� �ވ����V>i��W�t��'3��`%Fd��̞~i�`Ӱ��a�E6T�j��4�<,H��nx�����F�E>#CˠuJ+�`"��4.�K��g{G䬊s&���be��ZC�g���&�|'˻ ����'�F�S8�z�"��,�6p��w��\q8o�C'�/���J��[3  �BqG�M�������-�y�7p]	0���p��"�ٻ}�/xK�@��X*�[�����'2p":���a5��o���k;�ҽ :ME�J�&�����2U���<�z�l����wAr<eo$JG.����E�fg��:Z����Iu!�1I��CMt���5"/�K��kT5((!�r�(V��$�X���aL^Í�3�},�+Ǒz��*-��f[;�KT�c�v�/C	�~i`� �WF����A7�K�c�{���g�a�����/[k��jO8\߯��q�h��e��eÄ�`�)D�6���L��n�o�f�m͗i�ͅ�Ww�V��}� �/dGp�z9���u���s%x8{�m=�\;��I��n;���=qlX]�
,�����p��2����r*AO�j0�s�
2��l��W�	Fڙ��}jTͱ����*�N��:��IȂ�Q��[T<��Y
����[;	�ˈ�xM�������Xf�;��1|�����y���*�#x�I��9����J�8��wV�,�Ų����`}^�#T�a�s���9{8��}c�s��w�~�g;3��`ŀ���K��z��1A{���<Ɲja��V�A0��9�?u��z���|�<�R2P�	�,�Ȉ?��<c���KY?ӻx�U���I�n��^Ҽ� �ߴ��'zޖ���7���*0�/�_���<�^R��t��5��E.ӤR��^�p� ����
ϗ�թ��@I2���Rfe��'�Ҽ4�Wx6�HL�k}�&�ԙ�5��&����G�����T�
�N�ɜ�����;z�Ya`춐�b�h��o����eЬs%->ׇx2���J�E� ���%��f��	]K6-��G�N'���e��m<_B�.�9o)�5�Fv�N"
���BC$y�{�}���� |�1�3c{��_�X�)CXt������&���2˪ �p�L����yj($<1c�U�<[�E�dC��RK��AG�++���xU��1��M^|]��iH|�+1�.=�sb�������*:~��v�i�Dv�류��u3�d7�-�hW��5�"�ct�����`�!����������L3i��"?�U���]w�}f��u�F�~���&?���p�e&NMu��Tz`w�k��G�6ꋛ��Y���Ӵ֪��99&X"�@6oQЗ��R�~y�J]���&�!�A!ܡ�;�|>�j�-��	����|�b�����[�D�͙ɔ�lV@Cύ�)�G��u���H�2���=���z�NKi�J��J����u�(�q�p^Ab���iX+7a����9�FM�:x�^yQ��tS����/�⤬ޫP$�b3�S�;�G���G�_��j���4iKk0�n�f�:+�R��fP^��N�I���T`!y�a�	5 �ENs�ʏ���i7N�=�B���	-%�	�$$]�c��Dۿj�.T���t�]BW�E	P��N.}�c3��RW�\C&�D1���\�;�_�&?t(Nv���������_� h��ɠ#a��m8���<�����H�nr6KKy=6�#�0P�	���������]�Z�X(F>���k(C��{�3�eC���xL="�5��hQz��o�]h�U�"{G�#�����0�J�Sl&�ZΐàE����L��`g���sy�J��� ��;�u��RY��~��v�'����>|�8�\���~�ԥ����=�9�0L��p�@F��Ġ��7c�����uel��Z�}�=L���S�<7���}Rz��#R	?���2������:z:�h�9�7�ZBc����J%9���`AgԎrwܮ�M8ܓ�>�Օ����u�W�G~uMp��u�������G�>J�����ʎ�i��׏�>���,OŞH:��y~�nR��0^��9)eN��k�QhA�@��m������22��8������vG�,x�˘A���65��0�q.*p��V:���d��q����D��sJ��ɚc(Ry��j'&���Q5|�����B��ݫB5Er��J���=���x��92}�UXIFn��X��ap��.�
H�eLQ��l�