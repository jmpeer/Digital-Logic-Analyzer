XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Hn��[☫dZ�\-*6�c�=�(�E�<;�~š�3��S�K��T~{�j?g�I�nj_s��cc%�dEt���wL�A>4T��L탋+�����qY��X�gk&�1�:�؋^�=�Ц}��S&��@k��/o��L��0V�O6��!���!���?�%�@�F�0gp�|L�t�i���`J��_��jm��Y�~u�Xt�b�@M�:ė�ۨ��9i	LN4��#�v_�5(H�����~�ÈM�r{������4�`V�ac���`T'=�N�)kO�c��ۥ��g�`ދyC�Ўܚ����D�׷|>S��Ł�3�+�ѥ+���i�<�B���woW��H̲���h6��`���������6s|�`�p�~�ϏK�P�"��ts	a��$���{~���L<�F�N3{�Ўe��)ҡfd�0���p�f��VUWI�����ڬ?��+���G�g#�_�	����3L,�}S��=7(Q�Q/t�B�S�߶U�Wy��[�~|��9��'��`�
�c���_����3�c4��<'�QaM;3"�h4ξ]%w���Y,�H�@��g4�0w)\(��=���vX�#)l���zy �|�O ���J�N��!a�?Fs�l\ob,�'f��:&�1Sk�ٷY?蠉YC#��L�'��۳���o@���U'hj���g��7�ϒ��O����CdV�}<�i���P��j��3A�G󐰫F�B�mZ�_|��	��XlxVHYEB    56d2    12a0Q��3��ƪ\>�r�#u�p� i��oF��D3�B#'!�3�3����.5��֨�L!@(@x�@�ŶC�ӈ����si֪�(���qJN�Y�I�Ö2I�	'�b;�nތ�j��T��Ai�'+�)��U����y�J�6e��d��DO���&�������0S`�$g �J=`^R|��.�}��I��z˴�/�{�Uz��ofNt��	H�O���ŏc ��`��c��'�z-���~�e��'���i�ob�X�Q/�55�R�^mأM��^�jB�����o�Gl.�0�lE�R�#�q�Xa�.�* ��8�G�[�d����z�:{߽Il�1�>�f1(�[:0<����<AŶ+I��~��s<��N8ץ�SM�[Q�,�z�E&�haKy�AA����OSw� U�`�����aJ��V��T���n!�	X&�&���c�W}B��{Ns)1���yӑR������ŀN0{ȇ��јu��`�HU���Yo	,6wZDA|_;�����GI|������Q0Uv�q~�๲�h��l�+�k�Ws-�ߎ��s�������F�'b@����cmp5��h�Ѕ��I	�O���;r�|�%���-K�=A��o:���{qNhi�i8�7��_�|ыjH�9]����`����������%'��<�o��ifG�U.�I����}u��{���L�a���0dͰ�(�,PT���+R���#��VJ~�9g=Qz���v��eo;�)�q	9d�����08̏�0j�\��0rX��,��Ť�G]�� 8��~���]�JZH�� �1"a��|&��p:2�4I��H�.�A�T$!����F��2�;7nA`	s5&s�,��I�����z���Kհ+-d#��[�h�	 ���k�@�9�#��	+7=;uP3�yN��HH ����^��1�?��R�L���Ҟ��dn4;�Q�ઑ8�,�(8?�hg���ӝR0`��+._w/���1�>}��֏�`Xx��ox����)�!߸?Z�Y;�/��1���N����o[laK"'��lGٙVAj��A�O��Pz��܉e<B��'��v$�5�6����(ٺ�)'�����ú��& ��TP����[�֙*�{��'M�+d86��P��Q�C�f�q�S9K�o@��[�5l8ѥ4�� ��,����<��<.R0� �ۦ��ǐ��F�Y�Ez����A3��4@|�C�z}�^�(%�ET�5k�o{��}�|&ؽ�d��T~��VnG6��?AI���-zE�\ �*�|	�9ʻ�MK�5�Q!��V�[�?bGʳ��#�N�$H o��M��x�{�n���m#����c*V����?Vvȹ>.��3cbd�(�����B�/�(�,�����h$,]
E-�ϱo�	�b1�\p�)�
ݰ�!t<0� ��+Vzo`qA}M�ݴ�:�ŉM�ϼ���	uʩ��x�k��b���7����1�.1����9'�F�$l�vS�U�9�Wj����2�7��vbO�*�Ļ�3=m�\����m�1���3CwܝI��P���{�Yt�-_��a��A[�� Tr�ռ4wM ?��z���"1˷���T]9�^���2��W�E6��S��c���7�.!���k̒R�B�VHѣAE��H��xy�:y0��k#���ڎ�-�:�G���
,5���2�MT�˝�<E&�L8����I���(<�o�	�v�N|o�x+V�}�.���D�Q7D�j����U��R��O;�4.������
��P�ےgݑdh�L~E �_J��ISt��s��3����5��ڨܗ�����O�`��A�z��!z�y�q�d�Ĉ�rw�J;�".�h_1JN{N[��wN,����fHlM�%~&Q񥯮3�����<%ySӎ�*����H$�RW5v�~�IT5�.���;s��P��i��mli�?.��Ê�4�HD���+zdԝ��X*=}!dK��Z�:���V�X�ǀf1�$Od@}�Z)w�yI�x���^����kr��^-�4�V��He�I^4��D[sMi℈,e��!�O��;��>��5��
H���[;G�=?v�%Z��%��@��~��o��&�d0�C��#��l��pބ4Y)���ލ9HA/e<-�M���uٙ?��\kH7$�d�_�������?e`#���1�lg�������S��w5S �]�Uf*��|��y���Ι�t��'�����t�/}[����&{c攈/^�@����8�>%��|�EG��=3�$�T2@��6�A��B�-X��G�i�M�Pw�[�9��� ٧��\FR�B��ϐ9oO����E̘{0py5g�d)�z^���vk���3�d�p�	�A��Qǟ�#HI(��x� ��n�M��/���hO�RMlik�����O�9�*:�b<�B�`�^���hY"�Z \�[�~��8��)#�	|������X6�ͳ��a����4P����?���HI,����:v.Z�\�=���&M*kS�u�WջL��: [V釮�a��07��,�����q�Oz�ci�<7�����E�*�|�����+$���w�z��\�����h�J�m=S\t�gŭA�5��R�����dP�S�k1�$O����"�&���(U*�I_;T5�����3�&�{u��a���|P5��O���)��qx�"��0��hm��n��o�f%���v}>��t��bnqA�FPj����}�=m�tZ��S%�RQ��r�������"��7,3�@w2��bܷ��JF�2���
^�Nq�r����������H����_�q�i��]U��5���)&2�R �[��W��iݼk.T"Y�~����L�=��	!��"̤������"��KC�k���l˕����tF ?d�@Mj�|�Mc��;��v�H5����h)*8'˫H��$��s՞S��1�u��_+�l���8	ݠLm���Ў������D��$��AX���h���\sc3�$�[�s��^+�D;2�p��7Z-�#f4*���2!q�Aƴ�<w�@[Wʯ�����QZBb;/�E�P�$��4���"�Mi��?��Q�5:J2�%��xJ9w����)n�o|Z}���`i����������<W���r��kaD	|���W^:x�K�*Ah��^��k�|@�Es���a<���t�S�G�nֽc���բRs�YR��(���!	�`�"Ll�?�v-�����ybE�6"\��o���C�<��Jj�rs+zl-v\;��5��"+zdP�@�U&co�b�,.���:b����ڝ~����;gv=�A~
k��=9R�-Y(��g�qO�� )����b_�#A��_���Y�=�/5]e�a��~3��8M�'8�4�p����t�px�]t�?P��er�	z[����>��Ma�_!�I���ժ���V�2)b�k)F�h��G����+���}Џ����Z=1�=2�W�5͸Op*�x��!�ѽ�c�`��Ρ~�-���/'��Ǡ,*KV�����Η���&�km�H�D��҅�p��`hC��nͶ��nM$��!(Q�L���b���U�ׂBz3�J@S��Ï{��v�9��m�{�����c��};sO6+�q�bI>�iP��Z����u��_д�ך�@(�6X��u�B�3�+��?�J�A�-)��6Ϟ�Q�g���[�1NQR@H��gz>�D��n��	��l��N ��M�<#��I��Y��u�^�Ѡヺi)Xѹ� =T.9*3���ٗ���#״��>�)�-3~�� ���['7	Z�jO�b6���^�\a��>Ul�l����<~FC?p9R�z��r꤂%�S^�����x��K]W��\���J�QQ3/�li6���b��%Qŀ������"^>6}��G�۶:���b�Y����}y�لjO�O�y��[ѐ���u]yM�z=�yu�5�]_)]��������~Q��ؙ6z�����/́���ʣa1���ǖ��W�{qbO|2��{��y9_�2�Lt�z~kv�!��N�S@�1�;ӥj�N�37��_�5p����4�����*�u�Ή���
�ݎ�~�Uƫ�q�.��ö�$;��m2"7���o��`��&2���
���i���v������vf��)����L H�-�FC`�u�܃��+Ӿ>����	\�`i�x+Т&?��ma��r_<���*�M�17ކ���T{*+��u�^āV�n1��X���%�07�Wem�����G����BZ�Uor�M�ct,���6~�z��s8[�H��u�`~�}��7n[���ZG���Y���C�A�/嶼��p�8�w$
]�+�8��9��(Q�3����Ji�Rơ4|��Lh��
���X�l�Y��ɗ��KQ�rP/%'?W�'V\
�1��'�}���?�!�ZA�Thù>�s��,Ą,P�Ľo�4�E���(�T�έ�����������$�ס}=]5-���yF*� �q�8f���&�C� ~��ՠ�W�w����_͈�~L�Vf�c��;��1l��l`r��L�Y��TBܩ��]�����>G��:Z�����{���Qkڙ��ԣ�ܾ����X��U��2Cb�R�UT4��[~V�W����4����m