XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ͳ2�9�:գp7�TO�#J˒)�/G�����׆�j�Ѫ�V
^�����X�ur4�̠���>�eE��I��`��_�C`��?͎�@ FB��9C��ST�M�Yd��aszD3���^)���i��(
�����f��j� �8��MG3'��	�S�.����;}֘4���j5�aI?�����c�`��At��Vi[�_�B���rph�B� ���_5�Rdn�=r�� ]I
0M��T����ym���lk�r�o��W�-��=��s�yi�Y:Օ����q�讙!��� �a�<��]6J�֣��-ԏ́Eэ�/��ڌ�"^"�RV���?P��Ƚ%=m"��n�����>��Hd1����*�3K�q�IEv̓�6�~�x�t6r%Jw����U���v>�ib�|��eZqN	���r�i+�#��u��[@ΊI����T���2	���W��d�J�3��!@���f�v�
P�oY�Wcu@�c�˭B����}���	&��7����0�����obz[���,+m#��b�~�/�#p��#���<"M�q,�@\$/~٩�V�,B�F�2�|g���_��a��{�"��
��y"z��e"
Y"�����hU��S�QZ�S#�P�kYܬ�,^���vPl���{G0�՜���)��X��G�rj1D��6,	���(hr�����SQ�7Պ�?"̠qXRr :�6��겁ڙ1Шh�꤭Z=#�T�Z�Z�&ft6XlxVHYEB    c3e8    1d20t�Y����f�H܊5��
I$�(q�&F|�\�z�9 �W�>�Q�8P���ihp�۷+�b���'��}y���?�3<�H��Ub]�pK-�u�E��H��
�݌� �7D����L�.��V�t +�±=�f���R�g���g��C��O~�J��Ékb!�n�Y���ب�h�	�F�(΋�i�=���TO����	/���ɖh,Oi}*�-�)S��^R�vY,)����
c�\��WB���%l��;���(:��%PAP#q��fN�z3�$���\�#�L��,�����W ���~!��@�.5A�ܞ� *�n�AɌn|p�류zOL�\�L��Wl�ű�����s7�~D�u��(��A��GN3�w�)w[(�=��������%&��Y�i�H�kR���T�u�R�`��I,U���������4�Ix�nv:5�"Z�m'Q+N�}a^�?!��?vl�7h�mI��^ޏ'{1�h��R�M.��L�P�����ssm�L)ِ�W@W��BX����x��z��	Ae��de�Zj�r�q�OF�;e%e��{;}.w���`�3���wy*��-��(e��O����V�y�	���@�MX�'�/�9��[�Q�<�]A����4f�UN�`�$1o'�Ѳ��&%�~�R�O��MW?Եn�Ձ��~��u�@&�������^x�A��ȄO7�W��΁*}�k��[��;sBن�B�̾���hCy����Z�Bb~Bx�P�*L��`,+�H��OuN��K]��#�
Jo<&F�������%���k	�T���!A�-��@��{�Y�Z7�����ע j��Y����{�M�����G�c�,����O�`t%Q�y)$�]�� XI���ֿ��ڲXk����˧�J��h�["�x���e��Đ;�f�䮭��*M[�x��ZreIEA+m2���7^�xh���C;t��y��h��PB���#.����w�ٸ�IX�#U��H�_Kt�vc8�3�US�TuB� �7������� P.�YK[5�A�!ҟc5;������A�Kʭ���v+��B��RUzz��H��X۷H���6,�Mdp�upZ��ܷm�fj�z�ZY��آ�{�R�R�/]Wk����Ǵ� �
{a+���GD���ju���P�}������"p�m�L��`�^�b:���9�g&f�^�k�"��3�LeAJ�L�^�Cܮ��x���+��t��L1d��*�!WM376���Cswu m���,Z�Eu��$ D�k�m��㞥X�i�y�}�n5P�-����U�`+~��u$@	�ڼ����1Ceec_F΄̣�˖fh�,ԓ���G��D�)
�\#���Q,�A��f|4*{-K�nOG���vcI6W ���u$`��j?�d/�K���|�H�����y�GpW�WY�6�tD�FrJ����%)�	l�px��	M��nQ�d��P���xPޔL�f�N�cܸ)zzh`:I��w7����ة� s>�R��(7�����˂%�Ś�S�����&��gT�FE#�\�f,�hf���������㊷۰�b��Yǿ|BHRh̎E��&M���%y�#�V���Ï�p�;Y��pB9��Ot���5�a>�/�@iZ
�3rF0e������I)$2M��~�:Z�߿��ObmaE ܗ2��ɱ��,2�걮=�`��޽�� &/���hH�7��ꨆd�x��� #�$���(Kj�6X���el�9�U�]��[M*��{ÿ�ZʼW �n
ׇ����#TgO�E���f{�.āh[c�R}��D@�aP3CQ��T��{y�K,NU{����h���Xy��F�x
�0	��OC�5L�7yi$�!����/'���(������<C�sY���@�U�Vw1���S�����I5\9A�7y�@w97pA��x��Ǖ0g�I����@,� �&�v��G ��{ql�9�ďi�f'4;�j���ĹZ�t~��C�����������9��()�׊ͨ�QV�DKM�`;�^�ݥc��b�ou~�7��k�mtV퀵�5zF����K>��u�>g�e��ۯ���	�w��pX�C�?<���	iJ��T�֕�b{f�9W�xRǼ6�1���0���Qu�/DQ�]5������I*�_�W����)YY|�QX| �/�]jЪ���ah�ƯK1F\��'�� �D��w�r�-��c�k�l51;8jj����M^��
<���eh.E�����)�V�P�8Z�s��ed���� �u�!�u����
id^�p"j�z��.�F����{�,cX1�=�?3��_@�w�RJ��$g�j*��R�����s���`���3�	��/�Ă.\�%���ױ��~9a���n�L�[��(H�9����٬����K�2@����]�"s��XK��u��C:�{�e�p��k�����o�L6�͏�d��n����f�W���*$���`"��ʩI��(��J�E>@/k��ൽ�a��.���	R�b�J���Y��Xb�!����9n�|�Ï��s:;�m����
��j[_)(�ƻ��x�ک������-&2���2��!���?!�>��a�[g>���|�Dj��Ij��&����ȡy�X���-[=�0҇'��(i����/8Hs�hgG�j6�@��f"} +Q�)W1 8�eHD����L�C1I�M?��>^e^D]�ԏ&X�v�U��q���E��/R��B����� +���k��v�rΛa a�!���a��5���Qɒ����<X�]�lg��%�7�pg�6�:��U#E+E�P����-6�$���ܭ�|;��YQ�J�q�������՘��K�O�Y�ٯl�#��y_�_�y����� ����C�!Ձ-���_i��{
V�+�'E�o� ^��.7�7�y[�i���c2\V�.U'�9࿣���"K��i�q�gg���]4	��r栋;J�CSLD^%d�PTٰR!Lw���0�g�.�Ғwś�.����>����t['�N��By��Ska���L9`"�t>�q����2x�X�Ȟj�8s���Z�g.�����=L8�.�{<��;�ro�?~�ZX��`�
sy����%�R�F��`��5e��]�e5%�����h��[O��Fu����'O�u7�ڄ �I��ߎ���>R=Yd�X-�0*|�3n���NtMZ9�:�|�(��.6� 2_��(�� o;��	��۩k@�D���l�4�p�:v�cno�D毁Z�bA#D��ۜ5�j��q���YB�������u���-�@�p�x��l��d o�ydŷ�k㥹Dp���;�`�"����L6��HS�ոa�Zi��=�.��a��)N�X���p)w�y��i�}��1���?��(����DXQ�E���d[`��{]u��X�s'�����\�1>pΰ~\��DRa�/k�����e9��`*�?(v́O47y~	�k�ꦼ�X�A�k� �jZ��?��Þw�o��X��chf����{���!��H����qǿ$����/��7�n|���W���oe
��_���� D84*YHds{|.;[A7�Vx�=i�Vc9��Djr%��EwM��q�@�t
���,��#�V i���\^y�T�ƴw�\�]�N�7Z-5椎�-�x)0�E�Σ�R�Г��N�����a��O��2\���9��L�͸^o-�7;��9�{�$J�J(j���#�c�2�8��Ys�.���r>��8/!�fjd�f�!.���ʦ�̕e.���* p�׫����!y��2&mTu����^���S	�������QV��X��jx8��1��ʟv(?�S:#lh�d�ϴ��
D45�f^d��V3�'�E������l��5l�{�܃ۛч��9�8���2#{{����,���|g�����ՒW]e��TO���J��>ߺT���|�-3K�.�;>�֏\1�&���=���C�k$�&|�9e4���[��y���޲�iHݺ��2P�*^ϲAq�Fizyx����4��\��N�n_Oo��@K�g	����1��3�
?����D*�w��D�Ob�&d�i���w�&�����d�ժ���X�4#z�{�G_�Q���ɸȀSPp�OK��ĥr�rj��j="#�>fpb6]|^�l����%�*D�xq{��R7�͝��xbY4�Y��ވ�Ge=�N��T��b�`�T���P���.�)
��h?�V7�|���叆ͫ�;_YOR�JͅY-NQ�@�HfѕNYO�%��Sq��fm�ί`��UdL����zپ� �us^\����{ˈϡ�\(֬܅v��I*�2�BX(��RVIw�Ɯv<�������0u&�t�nJ�=�����z*p��,�9��{lv'�#Nө�B��`?����ɤL�Mb��������!a��]��Ɂ��9u�L��G��vp���;3J��8��
mb9��m�A�ӿ��+	�s�9����<e���\3���\
���N��\��a�� ��7���0�ym�|u�u�����h�l*�/�w��;������*�E���b��N�.�����Z>�b?�Vpk.��\���b8m���ֶN���.��	5�6���w�����z���e9<l:o��9�i�����He��}XO�G]?C{5�W����'�������zt#�ցK.Ϲ�M�|j�}�j%��1���G�
Z������V�����b2�3���P�<��L,��ǣ����@�?2*��4�WE^����
`>n�Ħ��FJx`b$��j3�f>�6ڨ�:ָ�-f�1!���h
�F͊�N�40z�9�7Bd-����.�`P�ؾ�Y(������wʣd%S'��"ċ���Jy�9j�q�ڶ׼h�nh_�q��ɱ��l�7-~��#��@T�k�8����5�J'���:�`�!�B��	*���ܸ��{i��k��-Hm	qF��\~=̒m��<����TY �oĩI���,N���)f�Uu/����h�`u�.�Q2��q{S��P�H
뺛h��Ł�zο36�	�lt]ƴtd���Pty����S��(IW�4�R,}������[]
~���t�.�b
�����]�I�LDP�Nz ��#z��
�P���k�&���6�Mٱ%z�(e�&�0��q�i�@gפm]v�e�N�JҦ�T����4~7��U����X����Y	%zZ��n(�ebL���P����<M���QDo?s7��L�\>呺�8��9}|ufn�hg�� �u��UAO�1��C3���a��j:�b&�v(�	�(���r�����U�Dxԍ#�TP�0S	�eF��'�\�͇��Ow*@FF�d�G���X���x8{frOA�NG[0l,���wQM�B{�z�$m�8�0��(͝�6���S0#=��4��J\cA���?��W�"����l�Є�Uq��v�χ�%��V�B*�L�kQu�!<�����1+w������p���ftcc�)��Q`�n���h��m��Zdު"2[5e2،ϝ�������˅}Hfq��l&vCƎ�V�da�wq5%����҂�0��Y0�?��b�K��E��{��?N.���J�KE@���(��[v���R �/3Jϧ(�$���T�$�_�^�7�����:Ip�!���u�ɪ{�4/�	����r�e�^�Z�:�zc\	|qG��ߵ����.�������6[���ku
p��@�̼W׀��s"%��+f����i�+ˑ��ܣT ?r#��IT@�}��w�V�˧���"2_��C���׬�JQ��3衹��%3.�F��ԌBzuu�3���������˄�Q�C��)�9q1,���-��ym��X�UK�s>f2+M�8��[-�
׵K� ^�G�aj&RD!��@�Nh������	�hf�x��P���&�����E�;���Ֆ�v\�-��н������=�>�pK�G ��5�b��ft4����"c	e�[^������><ZJ4��V�P���f�H�Xkb�o�>�I��n��������q7p9Z{!w�ܩD�ZᎳ�j�$5f#��u�0��>�P��.�X��d��]�lj8�RЛ#Z֔w��?��]���eኜy)A�u�?�h��a��A{ZZ�q3��GR9��W¹������!J8iRL�7FF��"y��a�*t�w���qYnlx���ѡ�������-7�n"\��..gÑ�j�����,�_P��2yf�u���0���n��*�8Ʌ��fTش$*�Φ�..�����Q�r!�i�;&޵i߯��o�B��	�ϙ&����srM������,&��8s����^�]Χ�8C|T��Ki�_ޢM��u��X��cTV�HJ��5b�bJ�|�oހrL�������j���D�� ~�h3�cp�L<� F���k_�1���4!"xb�Q�]��|\܀��/|��j�*+ >�W�Ĩ�z89{��$QH��7��J��:g�g�l�aW�e{�"!��0cBp���>���B	0�f �|#2�%tt/�e��D ��Χq�˥�mC��G�6� c��6�k}1�w)� �w_S<�y�?��8F�[��""f�����!$P�7���׶��_^l��U��F��洪r7.t���3��gVW>��^>�+<�&%x��iz�Gup|�2d�0��۝z,��a^�f1���Z��_
D�Sh6��	Zu�}hk�N�E\��{2> �+mΫU���J"��c��;���3t�&��4N�p��}��"�$�-��?T�-aF��y��<�K����k�ຠ����)@�[[N3��@�{����c���Ǡ��NX���@��=Uw�����`�Ɉ%��t:�������
z�]���%U�o����9��������W����<�kdT�U��I[t[~W}{G�*�_��t���U�+A�,���aL��i��B���fq�/�*H��|���P"�mM�=\�S��XDBB3i읢�[���P�s���m��v��=f'�	ɲT�>���˷<� �HO��N��^_kE�8V�6Xf��EKr��fl �o̪��+y�e��U��OJ'��E�hqQ���7���n��(��/\�E,޳.�a
�3_Q<Q�5��<��v2�_�9����H�!6�j���L�f�o��J�8�q����;gŠ�r���C3n��V_�d��5Ώ�j
;�qըS\�A�*YW�tF`�`