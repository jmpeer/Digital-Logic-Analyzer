XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ƀ�՞�������?iA�:�j�Ep�qPZs�%*L�	�H�E�F��|H�/P[�i�צ����s]�?غ�aCM3o������;�4u�[��8FL�]��۸�Zj�w D�qa�~����&��McH��d�0�#5�*-��u�נBLw��)��58g')�����sK=��Y��ZC����Y��І'�Cn��6)Þ,��:���X��o=�i�ּ���ۜ���}�̐� *@$���DuK;�R�;hf��C�
E���m\�w��n|��do�'j�	�V�!52��S�j=��x����lw��G7�m佬z']mo�nd`^��وRһh����\șV"_r�z�m�	�Z�2%G�sŜG��M�nQ���׃$z�����#߀�ʚ�!Y�ak��|*gCD����9u�)ؘ���quE�?3w��F���a�
ߚ3,�=UK¡��
5��,X�3�4[��W�f$>��ud�y�)[nYE���m�'#����p)�K�N8k�X�=R��Ñ�5f1z��a�����/�#�o�����W8Y����]M��ԅ ����(O�[zU���'�T\G�C�-ĭX����%�}�2�s(�#t�8H�^������8�@:��h$�9.5Â60̰��vs�`П[��5�{)��u�o|<3�x��E���l�����c��n�e�C��5"���!"���w�}|��cֿ1+c:���BO3S�n{��e�D�w���uyɍ:�D=XlxVHYEB    fa00    17901�J눍LQw�Q��9�s\wp��:��ƆtA�Ν�゙$@,�r���a�81A�v�����7u�q:/H�� M^Y�8�B���i�\�J��ۇA��o�h|1T�Ů����#�ss��W����B�rYۆA�c�kp?=�_.9G��Po�����Y�]gh�Z砯���v�@u��+&��ݍ�-��MKx��"<d��Z�yzr��4���BD���Z�X8��t�H7�٠�b�*�����%�hV��#.ѿ�y�"�gG�`��/>�7ag^� ���AH4�6�����z��f(�*�>�ho+ߨ�����,x5Ȯ�Ŧu���>�kaH��,�%L 1r�R��Ɣ �df�Φ���Y��l�~	Y@_�gW-�
�'�UP�ۗ�jō�#k��o�`3i����|�X�6Kns�~���N����D��Ź5cb�[��N�{���e8	���,F$å?놬���elH(_�_!#��X����G�*���A��������x��֯�
?�}��co�����+�6�b�#�ظ� :ݵ��Z��CM�+v
�ampz�;�3����C�)�����e(�W&���d	B���s��`�����C�!�u�9��|����Z��Q�Y��z�����-%p�#~q�}�r�����Z?\�S�C�x*�+�/ɮ�T�z�Z!,����z5��*��3+Q��ny�?���P�ߏ�`�;�@��%���L��>����:��j�q�95����ǋ�ٟ.�/a�%�W7�j��%(��=��@�6_'���P��v�6���4�f�g�J�X�Z�\���X=^x�% ��%C��� ?��%��O僖�$Gt>_� ߘ@;6 �S["�@9	n�FMPD|�5�c2�%��,��$;R�)�^�x�!#^"S7��넦{��7H^(��]7T�$3S�nbRs$!�͑%=�3����m
�<�t��gkm��(qO�Qy:8(�B��^[T3?lD�ZQ���`�hO�,-8���3�_��~5Y!v��..�Ļ��5�s��aSMn�Ej\Z�l��&Se�W��؇~�I�A]ؔ =kVs�6��eF�D����U��!?������☨��xܛ �n� �Y�!�l�P�=-�9�QXe��*��y`.����k������KH�t��#hu��!+��Ԏ�'0M����'��mͬ�0��n��3X�Tt�9�����˅��ZK�r�	���̄Q J�H_m��&j����K�aqqV#���N_I�?ϝ� _��"���iW�X8&�9���Q�����3���w`�dP�8�.F��Q����@�K���uK("q�ӘtuRh8=U��F�(���Юb�i�c^��T�+���؆��'����23�Xؓ{� {M���g`�lS"����Vh���RF���	q�&߹W�WX��0u���h�R�.���-�,|�5@�k���,��;�e.^��0�J���ó@�d<����se��/�%��� ��'9�D�6��/�..�Ti���W;�i<���P/�G��[]5!������������[�{, P�&���6���ԍ6�7����	�\�c���S�F2p5g��0��?o�@���Xx�̗.�Y�;�-��.d%�s �s�![Oi��^u��t�������	}��[ݥ���V�.c<:\Ň
�Ч�lv1�̐TI�'2b�/익N�ؑ�K����!5��w�E����S?Q@A_2�<��W�~z��G�_`1e��R?�Q/f�r(�k�Hev�0ՆI�ڱ�7g�H=�����_���m�ư
[�F�'W"�&A�H�qXWe[&ˀ+��{,8��E������R�sH$Jo[��fD��L�ǉC憛���K	Nb@�.l��Wz_�@m�^H�G0�Ȳ�>17�����qr�~��z��-����I�w�,B�>�0M����j�Bm_P-T�ۙ����fȥ�Џ)LC���#*�/\��h)9L��7��``���Ac~��SA�����U�sp���ۓ����'�;a�����A�}:��y��!����qǬ��7�<qnNį��ں���p�Dg0�ةy��5A�P��DK�BES?�#�[�h@�*=%�@ qO4;���Q���Ȣ���h�Ə�[޸ux˙�i+�&~턃�!�i@�K�!�W���_Q�97;��	"$����n��-�< �e��ɳ���	-�^�Dx��،m�&��uS�9y�Q>,�]K��Î��6.(�9(��z���ek�bn�!0
�4-r��x�J}���p��5	������HJ��7̪1��&/O%���h���w�[�0g�D@ ��)f�ҵ��I	�.�})����9��tw��Q����FO�x��O��eP�r�'D�:m�n
��V�՜���]۵��hV9Bh�(U�*�]a/�[h�L7�jr?ř���a�_���Eu�ΐ��D(�ߌ�;s@��h�|�������f�8���{9~�я�{����Y��e?lZ�� 
�2�������F*�	�;v�	�;Ǯ�Y~=��<��J��9��mG^�J����AЯ�ׄ[&��J*W:����/�T��&?O|�x��پ��I���{�w"�����!��s�P�/�[8�aY��L�7���0�]�����7в{:��6�j�TH���1d��[�b���嬁h�إ����7[^WM�栄Z�	��+L{�ή�0{���+���Ld6�F�-�ؿ��j��-��9�A4�C��U����� K��s	�B���e�`�����-�RF�i���C���.�s���Q%qP�;c�:Q(i-l[VB� ���	G6>`��Iú�F��Z9�<��˱��"Z#����Θ��?C-�*��EƴVͭ�~žVx5��^GBf�n��C&�2�p�(X]��i:ש4���&+Q���nVZ��'!u�0�HG�<]O���J0#�m@I3<H_�Y�5���&�A��a�:jˮ�O�/����:�h��h�i�ȅ�>���ʪUcV����_�Y��r\����)����rJI(F$����*m�Ob.�]��#�#rk�U��Uj�z<ԐD��q�[�f6��)�wx�f��غE&QZ,S�7���,ۤ��(`�}IM���4�ttXT�֦W;�������WT\����e��0��(Q���T��P#����7'���˟�`́�R/ߝV%��U��E��6�֌����b,9�~wp#��p����.ʜ/.�������>�RjR�!-_�@����r��`e�CiiRhaS��Uf(�6��#��c4����Ƽ:2�������9CZ]�_lV�.���ď1̃��������wԒ f�8��������_cy!���qݪ�o8�=�	 ����rg�{vaDl�W���;�H�t): ��?Ӯ�>��5+���
�5�o������3�U�n���;�9}��+���Ŋ-L��@�#/0��۷���g�@KX>��g{�@�77����B�"Ě�J)7 �E�w9gW��8SQ*���P��x��y�7��ne`� �WT�M�n�i>�a-ٕ[�L�G6�{�]%�F�8�Ig� .�!���I4f2d�=<]�x�(��<�Wz5K�G�bު��W
t6��N�$��x��r����"=fBRڏ�~����4��%�8"X7����=�R�7e��xu2�^��!g��'�Д����z��U��w���LH���<uDAx>[	ױ�K��X�[J���<�N*)D��d�>IVw�"���洆��fw�]�.�5i�O��U���"Кq/1a�ͧ�L;�&᱖g�/C1����ݼt���Cr��1탶�>|M⫶I���O�Z_}�H��'q�f�1t���:���������bˈ "8]���.��7ď����pnx�*�M�.�����o˹�}h1_�����7��/^�p��M��P�yۆ��g�=�&�z?�:��?�m�xr$�������=���by*(���x����DQo��P�:ę�!W�x�_�Y�|���J�ӛ�s�/�(}�wa�>˰�)�`/�Q�o܈��*ADu�|��Ƀ)�]^�BP�O�c� }�Ц99%D�a	���� ��p>��|����Fz���g�e5Ny%�Q� ��YϞ4A���f�Fۊ9�;�Ms� �2p�hs�*�����W�K+�����U�-.}�?����aF_�f1�5��d��T��H�{������W�F��o���B(^�l[��v�L۾:���.`�qN����}�Z������ftñ��1{ e0�����df�F�-�x�{&�LL�d5�{�x$����U�Ύˡ@�Y9 oز���\_n�_��܆c��J@���c�]��iw,^����]W�}��wP��f3`�]BTG?����G���3���	�y��o�);b.�/8U[�s`U��vʗ����MRT�s
� �x�Xg��C1�T��/D6?F��Qfn��Չ��6��4��m�e�~�g#%K���w4�!�#�җ]d9�nȰM�#�ќ��1<�D�?=�����_�zD�9�c_gA��h�S�s�
&vKw'$���y,�ߗh�D����D��{�s؃���GVekI,��Bj��������W�����TV��6��xa�p������ʇ���\�$���0�k:����r��.��������;�l��t�'��o��)���u���iJ���$��v1Ǜj"�l���XGK�[���q�+�����DQF��Lw��k�_��'�s?M�2�f��Y0��U.��i6%=)��fKr[Z :�K�\���I�vL;�rR��C�q�)A�x����S��G$�%�1��B�X�"L��,}�wa�`��R�d��Q���Ut�2�� ��cG@�_�pD���}�ɍ��-؝�	���˷SТJ ��>%j{�AHé|+X�"��'�fwK~��uf>=��2:�gs�ύ2�q�81��6oSp��ޮ~�p���ZvjT�> �����Ƀ���d� q��+p�iyXĄ��b��5�ك���G!L=���}��ε��C����7���� ! �r�"���t���+Gd�M<Xd��% �NUk�*�j1v�X��CU^��Ckٌ?kԿ���11N��7,�\K���7
�Ue�D���3�H�?qF��O�q�,������EgP�J�->ƭ@�}�Ir�J+�d�|ʷY���NY=
��(z��x��'��G�&9f̬J��P���!{�Ӟ>��^�q��QX���-��4|��nMvo7>""��]�P.����	ؠ$È�|�	ȑ��6�xb�'2�� ��*:��>Tfǿ�?Z��WQ���Vy�㯧�LI�;��s��	{��[�u�Ƴ�i��P��9�Xt_P�:���qI�,iwæ�1y������SQZ�ʗ�]|��!Cق�.�ב�8�ا����jdjG�*Р�X�_6����ϾD�s���	�]�i�f�;�A0q�8����D�EW�^٘]�fG�E2���jm�R����^�o�1ɝݔ|q=��n(��L�������;U��%P2�g�C=���{��~�|�Su�<�ji��r��g ��x`<�H����L�2�mj�B*R 3nً/ޙf-j�qL-[�l�%�QA��4��U1]�F��qk,�V;����>d�?�3���hL���6��x�<Ӊ[޳�*q?�����Ԥ��S�]�)�ADͤV��(d4-�n�(/ٚ� a=S��t�c�aw���&"���Ƈ����uuR��q��|�^��|A!��$_r����@C����c��$����e��y+�B]M�M)I��D���SQ��x�l��� cj:�����2@~%��ˁ�5�(��(p�zt��Ҭ����2_N��XlxVHYEB    fa00     5d0�D��^�eaT�pc��A^�T��o���}~D��bOW�c���*$ �^�[�n1�l&���9����`ϵ�]�� %н!v���@Pfၶ)q�K�Eb��t�nH�qM	�~�����U��r��;�̻L�1�K��?��0o�.v�'��<��4��{P$��R��w��M�6ف ����P���r�<y��+�h�a�_��ETrR��� R�����W��i�va��y����)�{�rr;Fy���C���(��Q=|^�΢I�_F�ƈ�+�oX�-}�I�3.9Æ^�S�nǫ��$+u�~m��}۩@���-�j�*d���фy��rW�Nr���E��,x���e�ŚF�)�����	MV��e'Hc��(`8ٮN��!53���6�-��p�`0;��Zk�>�ii]��^wbX!�}f�_/P1�?�:]o"a�mì)q���I����%��I�2ֹ�������1${3-���i�&:�f�:MUr�p���H��~4w���Z���}��3z�Z��#qm�Tg8�P	Ey���m�j����:�X��˟,^����X���GoD�fHoU����ڼ��ąS�]�YJ0�����£�lk��"����G���9�R[_����Dً���?�x[�<�ɘV�O�D��]��R`�N�S:>s�q ��1R�"8�=���b^}�9w�]P�cZ��7k�f�Ǥ�h��N��.4uWw���I#@: �[���W��Y��=5aFAjy�ً+E���_��a@	���k�ƈ���ԗ��$���EƎ��o@&<�l��<�e���-F
]*w����a��-����F]�������M��5>��r�Q]LrqR]��;�~�J`UFK�~�z����7�ݕz��E"���Cٙ�8b�;T��K�v��[c�F����~��Rp3��s;�x�ʌݵIR�;s�8m��� ;��z=?U���¯�X���6M�j�("TDGTWvht,�N����J����d�Ɵ����x_d�'$�{�ӫ�U��Z�f�i.�e��L� �����{����"pˉ#R�8�l�6��"�Ɣ(Y���2T�q&���Z��r	u��,�A���_̲c�:�T[{^a�H��O�5�g��t12���4>ۿU6��K%��k��u�9����e��c�=�nH���͊<�CB?�6�HS��Vj^mPtzzյ�n	��s
�����~A���klB�����'e��â7���������L����vF8{^�YP��_L�(Ϝ�C� 
B�ȹ[�]�7c��~ծ H5d�faJ��/S�0�f0����VVˆQ!'~_;H{�m��Sy|�>�@������es<za���!�j���/���}�ђr4����m9縫jm�ŮJ��#�NO�CP	襥�/LL�8|��f�+s���4����\"�BXIQ;yXlxVHYEB    fa00     640��7̃
U �>�W��N]f��E�]1/v�p2�Oط�}��"=lY�aQ��"�-
p7�y�BP%`2��R93ގ,�is9���-2�Z�� @J���kä	?������ue^I���̔O;$#%=I<F{�wϩӕ��-���@s��Qꓸ 	�V��@���Z��M~J��OVd���`U�f�����vF��-��B�
[��0�p�T�q%�����ю��-t�©]���v >&�۟�ѨWF1�BY�\���^o
�b�s*X�nK42�)�V�ܧ\����K���4�e\�D���g���µ;�����m��ԋ�j��	�q4h�]��� �3>�B�B�`�I�]&��cC������O�����1��`��Bsꦃ���~�;�t��7i\�vF�L���� f��GߊrJ�&d��z^ �E]gi抌D�$�j͵�PkD�oTbo���N���ìX6P�@i�T�"m�]�:�A~օUwe�%h�=F�6���Eo�E�r�-YE:l���|�e.)a�iU�wŖXRz'Ȍ�������c����� ��e�C�	!�..��Ҹ��:-SHS)��n?1��혡�w���h�yp���e�;�|DDV&V���h�&�:������F���RпF�p~ăTsk��I��ت�E��-�Kh�L�%����Z�����NBM�PVSM�P�ܣ�����H;d�0.��y����� �w8�t^�g��F�� �6��[@��w�3�2�n�:�	�	�$@Q@�o8ݯ�&� �G��\J7\��-�8JR
B���ش�=� ��(��6�g�.cĶ�,h��2���cvמ��ٖ��cϲ�u�v��� �V�0�+�|�]ɰ��f�La��/7���M��,Q�ȅ��5���!S�L�eU���J��e������!�M�YBj������ݬ�X*`�t�1�!-e�lC��C����(H��Z8Q��q�J�-���3y���b~>$-��8cQw�:L]LB@9��K۝�����m{k��cd�\�WErv#�8�i�RZ�dQ��x!����i�*���epT��g,�u�h�߫U�����<1���]�ܘ�����i�;�H����i�0�#I#w�t�6'0�Vs��O�%���z�H�!�sj���?�(�N=��};�&M[�������7��o�\�*<�^���É��]���Q���:�7�%Ш�i8�=M�D˼��$��'�3�n`��
헱������=R�*��)Fb�"�|�#&_��!��4h\��Ht�u�X#xr�����ͷJ��۲�l�j'=�q��vS�.P���0>�HL&�Y��iQ�x���ӣp
���b	���8ca[��},��W�F� "T}Z^'|�9���!"ď�<��F������wXK�&����^��$a쵠R�܇5�7�|g�5t��"Vc�}���w ���cPD3����Q��	O�jߔd#�_Oɀ����U�:	ƟVG%I�;������2��PS�`�@t%K�$�1d����%�`���p"�XlxVHYEB    fa00     5c0W��q����9F��q�=�P���gmH
�[E%�u����Q�<���ڝ$�57���>܊�h+��gXB�a.ܑO�7^�Ho��okTm�e\^\���Gf�	[nz�.�d�9�X�3�����H���e�����ٕKN��J���ԏJ�����ӌ��iQd����{�jБ2�H�0�i��h�a���*Y�p���)F5���P������e+6l�t{��z�YʝM�π|�&�2_+H^����-�WPh�1P�o^��+�̻w��0������
��-c��2kq�����v��9�MP��NB��k\P]o���/~�j���3E�K1��y2ຸ�����C'�����8w����X��~m22����d�,=
��Z�ݸ���G3�k��5Y��s�����T�t3��UM�fて����ͷ��������T0�����AW�R�
YT�K�=��jǒ���f?U��}�N�<hXoH����lc�-`Г#�-�#\m#�U�K�.�:���AV��W	щ��x9�D����X<z��_�1J�(��ש�-�����1�u �LQ;��P�
����WX�� Y�ʩ�D�ˌ�|�Aq��(j�6��Ė�ɐ8S9��3��G�?���� J�ɧ�>�D1d
Ỽ�Q�d%���Gqү=��+�A
������{���< �O��<�ك�6vu�Q�<��W�sFY����_}�iѭ�Xx�����5��/$�v��@�=�C�:I�Xj���a��`�sJiw�F��Ո�Ea�Xo*��I���K��x5���}�����.,P�d$�tJ�/���	��I[L4A�F�D��1�B<���.(��_�[�)0�x�"uN��)2����[� ����X��C	�V4���
�\,��9�tThpi��p�/��L�6(��96�
�H6r���S����uD��0%�B{2��=ဇŏ���#z��`�h�SV�W.O2M�Ϫ���^��C*j�ó�o�����bE=R��՛�K�[��Ğ�H^b���P#���1�pI�*:iq���,�~~�)�Q�F_Y9�׽��nI��z��U�	��6N�Vy��ρ�(n�L)r�͢8(n���|��������$.{��XZ�8�,���A~ɐiB:R�ʜ�l�gߘX�P�1���2��8� &��]�ѩ�Rl��2�:~bm)q .f�b^\a�Ix��C�=b��9�_��q�~:��;"N�U��k������\�:���Th�t�ܒ��kӎ���\�D'���s�PX��`E�Nr�ƨ4^�cu�!�B���j�UY�R5�^!ݿ�q�H^�x}-\�V�L�I�4�Г�b�4��m5�.iG�DR~���>2�qj�m�K��#�� {�`i�<S��������n�X&w��s7�;hg *{i�<�.�vJ��'�ؚ�t3t�XlxVHYEB    d347     a90��^1�`	�%X=�,ĸ>O� 7 ��\ �JI�K�5�eի H�p@�����5�}�B����zE�l�Ƥ�+���o���� \y��
p�/�,д���'�Z��G��E���H��E�V#����Ȅy�ŲO���bM؂�$x�M�`��;g��j�������F�D�m�/Ntz=,q�d�P�4y�6�C4|���@?K��҄FW@ћ3�2��<�%\�C7�h�zҵxd�1�����] �Ɨ/�ֿ�Wn���)�0��l��)��"�}r�	v�̏���։�7����jݨ�{��Pe�)��pe8 �'�gz wIɹ�f��ą���v�@��f�Z�:��2�;�jn���7���
TO@�[�?�N7��}e�SI��Lt
�&nvn��?4q2&&=��������7�;Cj5�r�w�\J��Q��q�\:�c#�T�ꆤ�F�=6g��s��f�BI���2JI�g���՘Dm�(��̞�w�l�[3����G#p��%xK�W�3U�S)�� hN��
-�xہ�00��-�X/��F��k֤U�v���O��@�o$W_B�8��x��ޯ��i�V�9Մ�q�>�N�*2�B��M�1P���G�j\�G��´�]x���f�\lU�P>C	��"�Wi�-:�Xq���A�I�/D\>b�Ni]b�`���e��Kt��ȡ�UN�2����[��#���t�m��F���|�,%V���[��TX�,�T1*��D^��5�N���-����z�H����T���ٮC���<+�%T[S����H��J-�����&�T���0�Э��������W��1�R��Eyȑ�k?�a�]�N!UU���|��|�<�m\l���W���b#zO?Z�:?�&����g�Tp6���6����m���݁%VI�d�1���ö��2,��?���%S8��P;���R�#����U�� _��D�k=P�ǥ���i*:�M�ےb(A���J�Cw��4�����&U�70N�YӸ[�t�|v�A����� ƶ�L.�G���^�Z���8��B��f����P^�Ƶ��5ށfh;�.�{���/����t*j�I9�#p=�bӉ���'B��DF�����/����r)Tz���X!@����w�K�Cq�����uWWp��'���IZ8fv�W���*��RK� �{�(P��+�=����i�L�&'[�\!��!�C��: �E⼰TLv�F"��K��R�-����~^���N= ��,�K�o_u5n�n%|r�-�Z��&�IL�q�`3TBx�(�ȡ��(+����B�p�s�<h�����3F�o�y�z�7]����)��Bώm'|y�J�b�lN����@��n|Lpm<R�����:ZA�o��Q�ǭo�u|�Զʷ�d��{��@�Ek�сBq��S=Ljg?_�%���͔���smCJy5�o=)�.ʜ����������Mý��گ0�΃���;m����4�ű��U~)��6���4E�u�FØ�)�t1��h]g�T=��ɐ��"�%�i�{#Md��D-qҢ��W^�_~�\������{|�.��#����'�<1[ق�A����C�������,x����.:pix����PF���38�_�Fu�	"Q옮�ڞ�����P� t�y�$C�_9�w8%�ˢ�˾�#�O^�(�Yՠ�B�o�i�"!I�SHq�?�	�g:�D`��D��,�/�͟X���0�����J�d�N6��9�+������= 5�����a�F>�DMOw#և| ������^^�;�m hm��zcǾI�����v����8@ZS:��@�Q�<i���o����Dȷ��.U8V,��Y�����s!���:�0��������^��4_�A�22��}�W_ks@�qޞ��|��¾�~S�cJ�Q'��'��:,���;��#$bћE���y�i  ����?/OPW*M�F{ �m#�TB���kG1���I��Cl���c�)������M�u�	�����HW^ݹQI�]�c� �brb<��N�^�i�O}�#����P��E��:��R�\��]-U��̈́k@Be2�ɠ�թ������i��3e�ԯY��0��|8
�!O*��ǮG̚��P���wV$CSo�R&�_�J����f�����wǟ��DuI�z�
�LW"���	���u5����DޖE⭻9�%tp���6��⏫I4�i�!�; �2���C��RE��:3S<M##�q��;ܹ�^��lfd�{�9;ڹ:,�WA$���W�N;��h���U�z��Owo�T�Od9��ə����%xi0�Փ�JA<����a��#��\���G!��T4�F�Ef��'���4*3m��i���������(���uS����}${���S�O�e|�חi�3����I��)Љ5��b�}�#�4H��K%��@�Vݟ�bM�h ���b�`��2\�� �mȜW���=���XJ���Y���8v� [�@��I��heoY�ՙ��m���#�Cz�/�딘��9���=����H�[[���$�·]@~�+��d�
O���^Vĝ��w�Ђ���k����l{