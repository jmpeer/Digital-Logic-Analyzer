XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����9��n,�*iޡ��M���&|۳�p~��N���"I��:���h��	�]Q�7��]H���q:�����+^��p^��qm:����;�w�� ��WjY�XE$�*H���6dO2��QVӌ/�9�9��զ��{ά���:dh����{���j-�y�އ��T-����o$!p�%��[%׸���8�ӟ�Ms)oF�z�)Nw��\��!p�[����]����b�[u���u��b�}^�G~�[l/0�{1Eb��/�D�]SS�ǳ)�{b3R0���ׂ���� ��uD�	�f��+򚒲裖g��fѻ�? ��5����9�6���۴v"��Y,߇�Uk,o�f�-)�Pg	���d<�B1�D�J�(/��Q}tht�3�ԧ=a�'(����}eKXj��G����j�;�]�S�C�)5M ;x�q N*=^&A��$�^HA*��������Y1"aK����L3�"ȯt�2���"�f��ex��Vm3��Wy����EQ͇���HC뤚��+=s�y��u@s��y���Q3�b�{�z�b���_ڔ��׋��=!V��i�yh�ޠ_���u��s�;;	���Aym��!��8_~2���;�";gS
�wc�ب꒍��n�qE��%�ޣOݭ�X}����Cb˫�\.�ꖀ3EN�p�6s��|��&��U�x4��߆:k���}�g��=4�햡ъbڧ�"O�7�Ӯܖ���S��&XlxVHYEB    4089     e40��J��UC�јu�bS@���{n��zW�$(�?'c46��&�ͻ�5��Ww.��e7UR^�\�	8��d\m_�� �]��{�x��X"2�zߜ���V&�®��VX�� �&������D���\3��L(g�y�Oc.W4�.��oa��5���C�P��C��q���u�cPV�,�����%���l�4&��a�w�����h�=�ԷHWT��'�D�lM�BJ��~�?f׵ ̀��5�EU��;��+p/�������aP�Wg�P!�Q�5�.0N��V-���kX�kZІ��/�䈍�j�Z�1-�-���<��]�y�8��r�u�S����{��p�vB}��c���]5���L��V?Z�/G��?����jO�H�^���)if��W�����1�HA�͛�K�c{r����ԥ�	
?�r�5|sȄ:�a�?1c��4�`DRή~i@��a��BXԼ����8pd��4���`��� h;�ȶ��m���OZ�d�:�T��uPV�$a'95(�E˄d�j��Y�����B������|}<f�9����z��"�z�|��B�T�V��d@�cM����陖,�<N�p�"X��BS��0���r5qwv{�.H���^�dU�Yd�0��@��'�#�8�f}���6��1?��F�F�|d,��
�$��A�ݝ�($�����zi����t� � �`�,���TcN����������}(q��5Q�x�S!�|�74Z�~���4e[���Ã���"2�pU
�߳,��9�~�t���/@�����	�c�3,;�	�%�v�t뢹�ܬ�2gz'0Կ۳zIFԬzX�Ϩ�PsI���y�c*k;��LZX�f(����0�0�G;˭8ߢ"���%n���
�t��,򰫫|�\����[:HRvOe����͙��ɮ�|D�K��t|n�����{Ͽ=�O ���.W�t��r�U�8.�6ED؉ �zqR恽u*�N�G���C\o�]^}5�q�O�\y���
i�B����h\c��rK���߁��/���h��ϪYK�Oq9�@�ݹX��҇�������`3`@�ߌ�~��?��?-_M��:���W̼�yi9�R-�4P��il��x���?~�9)� �_E�z���?ϩFxE�\Ͽ�K�� *�"�uQ�����y4ȗ��`���x��oQ��k؈�[�b��tsMZĴ���h*	~Xȉ+�єj�]�F�RS�fc��:?�*�c�겗�_>J��C�x(�ʞ�����?>���:��p=o�����qj���j��2�� &���Lݹ�+E�pBv%ubg�v� k;@����6����|2xe�����|jj/(��V�WCu�˱���5��.��`p]n��<���|tbQ��/_R���.��7�C�79I�w��q_�h{1n�׀2�f�EZ�q�"��HM��S�g��Q3pD[:ZG��÷C{<$+Vgb��^t�e6�� �4���B��%U��;��?�۪yg�K��}�*�n���`�w�nʩ4YA W
��@
�E}��V[�� 4ŗ���M��B78��Uܷ�96�v3�j�I����|!�	X�J�c+��{�hF}�=��XyU��5��{�a�0̌0����e\�vH�'�F��/�\�<�9N�����3m��uݺ�(�]��{< \�Ve�
\�\�*���Թ*��@�X��『<<Ed9�^�'V�
Q�ޠ��|��:V?�E\��,n�		�3�:?���-�dg[k��{D���wi��zt�A�W���Y��*�T{i��02���#�c��zt�ـ�p���?w����\�Z��7ߣ�K=��Y������_NR:��`%�f*(�]�<\x�?��?"!
�̱f�k��p�ŖC��*�W�X�\�f�,HP��s�;4�TOU��J�
]��6*�,f��mȆ7W�sN�&:F/�Q� d�aCN���劯t��
�USwZL5a����fI�6/� �1m�CY�p�5p�9�%�0�l�d��ܜvW�1���� ��8�Z�C��|}{ٯ���.	K���
��f?�qk�"�r����b�/����k}�e��R�{�����9D#��o�;l�ͅtٻ���ѡ ��f��X�;vX�o'�s� ~ͽ?��sn�TO���L��4��L�rS�w{3�aTB�$�TO�U2�R�m���)J�w����F�:)0D}�݃��.��)�[�HSУF�r�P�5���yTr�y�5�gN@e��r�N16v��S����%c����([��'GY��t
����u����`���'���yz?�ۮ�9�m����$���?��#gy�N�)��C���3жldr&ya���g�~~RF�����(��L�ٽx�k�Q>AĢÍ�1�A�{7�C�Cf=�$&e��5�X��{�5��.rJ>'g��8�h�T�>�pk��pr�Je���C�^*~�-���+�����2�����H�CB����Y��`� @`�R~�}��n�v)���^.49��p���Rs.l��0��Y�t�ՙ�17t�,�$]2%@�sRVz��EY@� {�.�� �uT�%\)�j�l
.▜��%Z�yJ&�i��P�N�r�����{�&M�GD=lhA�ǭ\Ә�=U�yo.�8��c���~�2I�.���Y�Ʈ�}֪^mM\�vDY�'��R`K	�Y/�ȭ���t��E�e��Zi"��){�IC>er�~p��UQ��	�Qj �[B'�mD���ó>����`�ć����[ۚ�jV,\����v���Q3sKߑ��`
�$E�BF���r��^���t��8!\ ����Q��al�h$�ٙ�R����nG0D��Id{�-xdv�r-�/m�?131�,J�ȾQ�=��-^�d��E�|�=�K5I�6�ͫU�[��4G��qD;��
�u ����'���R���#��	������z&��C�����.DҴ��!Ң��!ri��V1��.� ��sIT�qbu͌Tu����/I�U�x��,�����wG�_���"�7�_z	��j�QY��2*�W�þ�2̧T�\
@���h2=Z��n���J8���Bn,�vA=��;�N{�gT�X>�첌��@��]ބ:�=�����lp~�,o�QB��y[
]���Qy�����h,K�ޒ8`����t4��\D^�R� ��ca5a�]�}¸t1����Pp�ݢʟ�h���_/��UkDy�ǎ�d�q�n�gx�b%@���H������u�
w�`X�7`���h̐E�7�JPb�_K��=�i�ӈ;AGѩ��#�kH���K'8��d�Z�I���[����ImMd�'٢�ۧ<�9�y�����A��{�z�.�i���r��8��ok�L����֕�R;�Ւ�������N�d��$��ڭl['�S�|%G��N�^���4�C��jn�{<�]j��V�]Fjd>�)�ʞ!�c��ȿ�ρ��m�:�vy��P_e{����jv܄�U�GQ�m�8��~�
�