XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(�o������*�y� '�UP���%�x�$��={�@��~�������&��yF��4:����ϐ;�u,a��W�m61Zg�H����tP��Ͻ��g:�p1~�ܠ�زM����A���0&��ȶ��Zn}��
w���1Vg���/�{x�ߣ�[O�O��U4=	�8����3�D��ܕ�M�ʸ��m:�W�y˭Cфd�4f�����3!V!�5���F=5�iA'4�CA��U�ŹU��߽s�6���)���|�~ÿ��� I��V(����:���u�Lu��6 șh9ݺ��+�Ƽ#�<�iϻ���;�'��X55s�3��U��鵓7.�"[��V����a��2fB��Gl�r ����K�I$Jn��0��%�����,�w1�Y�������C��.�3��K��S�K�b"�k�.@,��!pB�@�&��T�[���\��As�`�s�͏�
_�{S퀜� ��b�P��eC�
���F���߇�)�_f��i�ƅ��0��A�"k���^�7Ik��0����V��HBX��>��bQk�
�;�B��H�ÀN-}|^3J{![������ɧa�Iɽ����3I�>QN$#(���I�@G�3ؒQ�ȤEJ����)��$4j����Mէ�����P��FX~���3�W$��#B�W��-]��;�IU)�\$��n8/�"��kWː[��/�tFk$ݢ�	�f��<c-���u,}5=�Y�XlxVHYEB    fa00    2560�0Țz�c�'���t��)�̱vP���Z_Đ����T`���ʚ"M�F�!׎4��U��۬4GB(�E.�-1�G��,�8\ k�c9Z����')��t9AHKF���n(kB��=�D=z?"��%fndQp<2���,����6�������(��hɱj�6SRϣe&J7IO<��0������KK(;���fI�l	s9�	�n��y�3Q�� ��V�
����Ov����"JCy��x�v��3��'2%��OF�hU	d7��*|s�Pu[��Q��U�ق�'��U��/9�m�I�l�-H���Vc�lP��Ei�����&�}ҿ|��̄���r��g#5*(.�������Eh�nV������d<bP{�̀�G�x`8���n@nw�a��*�Y���J��Fۼ��%`�qT#�F�����|�41���g�MƔ�t��u���[�A=�8������#~h;��'�F�2YT_�t�X^$�m�ML��0��� �-�S��Y꤫g��Ǆ�g�w)�SͶ�Ƞ	a�&�!�,�%�g]C�O"}��,��)f�M�
$�Ф����c��)Tɣs����_PI~j^����r�guNZ:�!Y��.u�,�4�y�����;G� R�D���Ǭ�dO����:f��k/�����̡��N�<y������.���&�9cM�I%J>�NSo��e��7O��`�B�V��B������(���P����~Z7&x�o�A���Ġ��;�z3�q3��ruo{d�n[�4}�x~�dL��_��
��K��dצ��?�_ݚ�e�1��4�#�����iOr=�����Ź�����t��y�� �*y�y���
�����!�ܻ�W<������-`BW��Z�;R�c$b-L�X;Z���'�-�����k�t)��/բ�	��it���nm�é���&�~\�CشEQ˿����^��~�c��y�iֲial�x	t�8ՌdGE�Tw�(�/I_�7�Vr�q�j^�DpV���c��k��K�����40
�R�����et��{:o� � �.�F�Twp*��]m���69�+㴋cmmP���9{u�)y� ����Z���|�����w{#%Ė%��� ��Vg|��ۡ�*�x�/#,4EŸ0p���I����,���Ũ���;���l���ZY���g��#�����,��]���]��Y�B�Կ�|dZ���r&�BB��D��	�%�g��C�3'
�Kq��̭T!��,"�8e����a_k�[)F�t��"�`tI��Y���g>9|�!�&����i!"|�R�	�Y��<lmF������Y9�&#�Y�j9��`�F���o �̚NzDH�=5\���cr�	Ќ��	��w�g�]<�Q6q�P86_kS������C�t}��ݠF3�gs���ПC^�� ��3�Jѐ�{��������7������}�i��a��p��ޏe������=�ꘪ!Cjʡ~$��h�W�yz����1$��>%[��Q��
FeS��D}$�Iݣ�6�H%�H0�P�+)����$��/97~t�&͎��]h-�AS�ZZ��i.������I�zB�����lR�:8�Y�v����~�)@B���7]$@�Y�������'�	��J�N�ڠ�d'ҋ�u�n�~���E�����'k����ON��# ��"	'6T#�~�L�|�I-G�S��Z�K]Mh��j%J|�Z2�m�n�+�ks�5�T�l�=�9�72�(���A�v���z g_�G�T�'���
Ag�"<�Vl�#DE��ɹ�'ʧO.hd�䋉�
~B @�D+?k���$�:Pu�?G,M��$sKR�E�YSc�j���P�:~d#+Hj�i��褊���7�Q3�MU������V�o�bń�,v��:��K=��8��k�����"���!6,����_9c��~���W=�D�a%	>~W'�'9�/�$u���G�')���T\���+R<y#=���QU�F��(LX�k��r����HȬ�3���@�<]�� ��N�F��s];X�;1�NJ��.��3�����;�5\�O9����a��:����.,�?�E�z��Z������పwڇ�6�@��q�w�e�=f�0�>S�"~΄Cv�"�v9I�Ī	�&�1mWw��������x^���vw�P����6�<A�����&��R��UG�Q#,��#�
��:���B�W�J*�C��0iů ��
��a��:��=�/��8�j�m��ƶw4�@w�u�����&GG:�E����b�X�sM�ľ��-�O�ګ�}��/�E��+�͝�`��s��s�ŷ���Ӥ����!U�l��sr5����im�?S"Q��?��ͅ(w~��לq# �?������+ېa!��-��k�3�C1�x7
��X�$�'�}�|h���m�f���)���Eˇ[	��ً���9T(�)
[Yd�pkb}�J��)w:�÷�����M�\�:�pW{o���$69�u>08��G�R�-����Q귡L{E}�
�PQ�G�D����Y�&��+{�gGm�pwpȣQ|	���_�ٴ{�To@��������
U=�yMb+W)�l0(�LBYLE4����b4mL(t����O��`�HҔ�i���"4-�l�K��
�`�`MQ�N��;?6�E8��A%߿���ƾ��.�����G��J!qW�ʍ~�Y#���ځg*�j�8K��̎SDey���%F��v�ҽD��R�0�ۍ�~r�U�ݫ���E��迈��/��PF8 �@����4�d��o��j&�1�����_�Syp�@$�և��[�Fy� ��!06�!��Z�ctA��{�yl�vO�/�Z�؛#�)��T����~^$����&7���l�Y4�~�8���%ŀ�q��k�]�<i&�&�3�h�-�:D)r��'��j�sf�nNk[�-�h�/#G�Oa���JR���e�	i3��r�tG���K��HW����=�#�Gj��y��L���9��v�pְ��z�]];�5/E�u('�1�R�}1`~^3OzX�<
'���%O��G8�g&ד��/�f ��L^��F�Xϕ
��e(�?�ۿ�*#�����5�c_��"r��"�x|��w�#Zk��4*9�n����,I�)�$�1���Fq�G繍�H(ܷ;�,k�L�w���=D9E	X����?���?���ӪN�u�`s1��Y�~��"ypPW[}>���z(~Ѓ1������N��"�d�4�Q�8x�]@��x��ϕz���ʸ�pD�fY)�{����Ag1M����Շ�"�d�L?��=�d��×%��h=L�l����t )Q ��G�kw�(��J�m�B��8���%WW�v�NK��K%��ON9w7�@���V�Q��B��~X 9�>-���G��98���Z����a4}^}��1��������j(C��52��5��~��qӕj&¹;^m������$Eb�>k[��b
���AL`�1tq��-�X���RN��r�jl-X�����W�C��� P���o���6R�z�[q�(=�ӻG��79>\!tFA����r8���M����TKlE!�Hw��9g.�uPx*�+b���_�F;B��@hW��
���_d7��p��U�����_"���n���F[*F(ֆ����Xm�J�T��[7�*9f���'wh�ہ�^�+��d3K�µ����n=\Q��[�!�K��HJ9w5qYLV�HF4�����E,\��؈������i!p{�2�c�-U5�`qHR�bx }Z�*��9R�2Ty0��cF�<��i��l�8m��EJ���6�BFH�ߋ91x�Cl���������!$e@G��r���SN����b���+ �a�/"�y���i�h]L�o�9B՛p�!k�M�[�l�~�{�{����Z.U,Q�BzNrkqٱG��
C!��t�W��Ǖ��e�+����f�3��`k�$'�l��_�h�E��>S�w:�2�o�Ax���;��.�9�E[=�T�XW�I�e�<>_�?���T���M�M��n	� ��H>��<��Q!��"�	���9ic9�H�f�轺1�t�p��'[�Yc���4�z~<z?�a�̳��S��<��g��C��%�>���r���V$�u�mނ���%ρ�DW�ɓ����Z���DE�3#�*��GO�z"��)��ڧR:�w}WWy?�V�$B�@d��ٲ�U�^���v���	n�Y��pK���_\Hw� A��O�{c��Ao]aag�����^��6捇���uQI�4�d��qQT��L�<
�+�����i6>���>�HF?(,��E��S��iV8U��]�.�w�Id�3A?���P���?�_����c�f5����iq�b,��h�צh���Ƣ:c���2P��s��4�}�h�Vb.��������<�̇�����JY�D�R6�e�ޡ����H�#h�j��x8x|�v�M��*r����L~��e���Ѹ��'*d��t��
���nƑZ�՚Ʃ"φ'J�>����?���9�@G(��ha�?P�.dat��I��K��/���U͇����9/��+���mn�� b�������Mh��f]���}�58���JI�p)�]�5�No�j@j���6{��%h�=��@P?ф"��"qϊ2�I����6���Yd��bl�LvKZ�ї�� 7o�p&V���:��f��#@c���,u�Y���$�X�<>�hDh���|���ŇdP�����p�Y8�eo�2d1NfE����-��۱��L�h��,�O���Դ����)[K�X)�������:=���v���<4���hwNֳ?�Gø�7�@@޺��>��m�Sm3?y~�/y51�#�c�f��v�m�h[�_�����C��X�!�w�h:�ի��E���,��>H��H�h!�����c�أ�b���K�+�g����p'��z'��e���zt}�s�%�2�/���E��Ҷ�� jp>mH�A-��@���Nc�>Ŝ�i�=�E~�M���#'?EίOZU����w����oU����Wb�0�}�(uR%M4Ȍ�RI�n>F[�e�!QcH��]�;��#!Sm�OB�f+�%K��{��]V�c�c�W�Q�e�}�?�5��ҙEr#�qߡ�8o��� �Z���!��2ּ9�+��C:jׁ{$C/��%b:��S�k\M��$�+��_gͧ��An�Ge�B���w�T�h���!Ћ&�{����Z�M�mZ���tZ�I�>���*�¹{�l�@�(��O���p�k3֟ߘ?1�z}$���?{[��Ŷ���-Ma���?�[�<�'�X�9B��7�AA"��'j�*���w�,D���ک���ҿ��x�5���Ov�j0DxZѥ��F���_����js\_�^+U�+g2�ʽG�o����l�N��cYL��m�k44��i����5N���FJ�o}���Bj�A7�$���L�b|z?�)1���v;F����H����s4��y����ȼ�#>.gBL���K�@V{��'���|�쪉����Lxp�����	�Q�s��vmĴ�D\�����B�l��ԭ)����mƚJ��Cº��\6ʻ���AR�H "�$���X��rޔc
"UQ�����`jG��A�QK��Ю��A������d�DY?J|U��%��H�n���HJk�g.c�myq]ϸ	���")��DJ�"�el�ԅ��IUb���6L��$�p���)��ߺ�k��"��M_zP�w�>�0A#���r\䳧7!�ħ&*H�P �U�=�/Ux��b��xɦ��-�A�:�;DI�d���bm�Ա�`�p_^���>g�YE\uR.,��G���*V��j�����}Y� ������^&�E��Y�<>��i_�M����SK`IA1�31�;y������@ �����{��PO�,��J��+��%�:�X ޒ���W��5��j6]��Ȫo����Ҟn�45ޱ����|�����;�?�ìX��;S*�OlR�p���V��q��ΎL�|d�#�FCe�]͖)��f���j|ͩ�/��#�3q�GlYl���z�g��X���mip�#��Ґ��` �J��n����4�v	ZwcY���-�n�X�������r�&NgS�%>x;��R��	�L|f�Ƣ��W��S���7�ڢt��3DǓt�=�0�v�L���O�bp���N�^�5��@�`���/q Q�S�Z8#���AB�*�9�CU"\$�Y�'�����[8P7�$qR����sÏ3�e�
��6��ʳ�bK4uH����ʛ�*����n��/ːI��!xcȗ�Q��\�	�k�@�[�=�x8�Irw<*yHbpg�X���R�C��3eӂ���t�M�<�5���y�����J41�J��#(Z����D������;t&&������1	7�^dz�}d����1}��q��0�k��hF�c�qΫl�ۨ���/	Ķ��~i�rn��n�z-][�kv^v�˹��-�֕� �t�e0��R���6,#�k�Y��&�ZS� ��P��,�5A2@�e,�f�Lc���ɿɆ��u�5�E�����	@��q��-Ē�<��&�Q ��俗�_�s7:Z���d�ge�b:�^��5�˨#�<�,��)y�S�.ZU?ݙ� w���˼]y<���RG����7�Zgf�yF�f&�&�s���]����(����#�rQE��J�En�����t��ٱ_]I��:��|Ъ�z43>=�r�%N[�kKO(�d�.a3��r�QΞ}4PË�NS�p��ygz�~��]�QD��u	�d������d����}+����O7{i�RSuIiֵ?�;���f�<�(���R|v������%��E`rO��d8Y~P��W�a�hZ��� ��}ӻ�Zk�����~�����p�s�[P��&�e�IR�ǒl(�c&����p^X��j�r�[�����iڇy/L=e<����c���P0�Aq#? ���m�b�b%`a��$@e���[0V����oj���E�`#l(����K9e��B�Ep�S-���E��1��}�K]TvM�K{�d�*U���ª���y_4_�äɦ��۴nM��@3XT�&�X[v�RM��ǐ�/k�ί�-�B�X%0�A���C"�Wڼ�;?���Wl��iu7�H��IM@���"+��a妣t��T��
$�' 4�j�-X@9u�srm��'��+b;P�>&z^ۖ�Y�}��:2y��N�����"I;�FǊ��B�=4Dc�C�b�U�T�b��p�[tX�J��*���,��������hRd�p�̙�+�geEؠ�P�{ll�L�W"�,�ٿ7�D���/�	�^�9��~�_N%.	W�t��DO2=~8���5L9�[�ߚ.5U$���)>m)�T��6w�>�M{�d߅i( ���ާ���q:�j�v8�9�@���Q�H��\�оaO�r_Dً%8��`����E�c+w�]�f�t�#��q��G^�j0Ys��GYA�ήi�L<˂��2�u��r�jHC�-�}��P�&!��BnB�_�+�'ɗ�qNʢ�_T1��2�;�OY9@%���~���K9��3.�A����DZ��kj{ǧ$P>�랏_���"X{Pa[�C�*�%��^1"�e2�b̉����r J�Wc+o����u�b��舾�j3"��/����\��҃D�Ƞ�����`�H<#*�~.L`�|o]�^���g�$�hs��tN&ᰜ�B2���=���+z2��R���[�a��x~�c���Yڅ��NLh���dN��:��{Q,8S�,+�Dm|�u?|��� �5Ο�Q���R����Ft�\�=%�H���YD��s��-�':����{۲}:���A�����v�-���!��?�R��Y��P�#�O��A�K��[Fi��0��_w{Q�6ŉx�����F���WG#~E���{�1:��#�-_����5�W޺Ɓ]"��]��0�S(�fh�[xa�xl2Ѧ���AC��:1k��#O~�zW��9*V+ԓHn��}�r�z~��.oK�*��0�s��&�����4�y<-��	d�c�s�RsȔ���X��i&!xl�K�Yt�\����(XKptZ���,�#j�O�0�w�ں"~�mҫ$��gz~����s8������:Z�K|e�>|tUԔ4<W����d����8��0%��r�G��q;/go4{{���0{>���R9��.�� �━
(@�����&�sq��,~�7O��o�ޖ�:�!X	uN7a.z��"��y��D#|Vh��{fNgl�Ŗ�N>zx�(]EL4J�o����dߦ	+NO1�C��]d�#-�l��Qb.�z�شV7BZ�¿�=%�H*x�u�����N4>��^؁�ly����r��b��ƃ���q($L�%�X(V�n��m����1�"���<3�-�Av��k`E�sk�Pz�Ş�$�����ijoW���I�.�F;lOM��e���p׿\����f��1�K��ʊ*f�I���ǵ�)]T��|�m3c��}����u�������Q�tf���Dœb^(���%�մG܎*�}Nڜ}\U�;�5{D���|�� �/����0��w���$����4݋6R޾�+Av�X`�fT$Tnԫ�ݎ͗�4B�O���v��W+��U�j�%�"�u��Ө�@K��C�r�x+yoZg����F>idM�ߖ�h��R�FF��ŵa���9��Z/2���$hJ�~>v��4ș0i�ȟ��o�ɽ���)�J�58��X	y]W�i�8d�GUA &�cOX�5�F$/A|K�Z�%�36?Â@|h�s5@��0B�	�;��(�Ѫ��N�����	��������-���뫲��j^�>8-��c�]�,%��!�WE���?�p� f��4��L�ʋ�u�B��A���'���#�K9����N9i$ɟ�Q���@�q���Vp��}�a���ȓ)�&�S1|�	Z�1�d��8p�y0�c�HHAK�����S���[m
�I�b��i�C�ď�X�i�E.�L�$��?'vT��:�o&00�0�Mz�R�?}f��L��xm��0x�?Z�)���\l�Z��i�S=̳�ylG>�∆��{�E���I��b��jQm�Ĵ�擵 nr����ox� �&3X�{���7~�C������(��@0*��r(����H{�iXlxVHYEB    fa00    14b0��!�䀉(��KM���~�'�� d�g�'�h$�J��e��Үb�K��M �o����5C��دy����"�̍W��dWM�3pE�Ѱ��0c����/�7�j���Z\^Μ�L�n0G��c��R���2������i;���;�W�fU��~�:U>0�;�*̴��W��U��u�.�c���"�������Y�V�&q7��!x�aB��$�b����Ze�ъ2�
��%�a|�'I
�/^b�Q����sm2�����<@��O�}��hYV�a��#{@*��	S��a�V�p���xj��l`�W��f��0O}��T
���=,�����������yYo�u�P�F�{(�IM����ܤ����j�b1/d 	�X�C
�+��c�RY�>n�ؚ`����=׻�F̷@'�\��,���"^�����?\D�?Ŷ.�<����e[��Pg��m	�ũ"qۤv��!��q=|qKFqd
irK�ua.�9�gY��x����4پ���e@��N�ι��W4�k�@�#aݗ��ru����ێԮ����*���7A�Ͽ�e��Ќ!�}M��:BE�C�"�A��H ����'[���P��GMR���5�1��X6`/��r��D7l9X�+�:/����Чz���WI?dK�`���qV��ZUC[G}E�͟8&�=�5��Z����g=ty���.sY[w,d0r��;(#�`���U1���v�p</���S ���m*��o���hE��.q��r]b��f�	�E\봰E�Ԟ<2�v��%�6���)�[J�0蔨V��Rt���Æ��F���C�D[�1R��k����_�i�=4,%Q+1ת/����Lp|S;���{��dW�v\�к��ԞS�$�0��thd^d��4cuK��}pك�R�Q��I��`O�]75�>!i��?/���T;=`�v�k;�~c���c�� K��:1Y�np���w2<�M�UPX��L�y�
��k�ݽ��/�ؒZĔ��M]u�k2����a��립���C_JG.����fhM}�Ԇd�g\OF�%�%w���/�������DQ�uo�9�/"���y���1R��(i��y� �(+�W�2\I�|Q�m�YfǨ��RKy����ǃ��4��9�vd˕0�s��&�(���i����SG�G���-�?o}����d���G%!�C��s�:���Y4�~������{��r<�VJ�R_�Q�WC+�#*pI5�`G��6G��eÐ����nzʔ�����Cғ�&s�������GT����S vT��oM^�~v����
�����D�G	�ic|q�r���y��`��Bf4�WZ�1��� F(�%9���Fb�����Xk9$���$��jj&-�n���6#��@�(6�|�p���|i�_.�5*;X�;îya{hxX��tQt��7!r '�"��r�&�����3W�#�yO0ͦ����I]�(�
����W��Vsj�#�_�]&&�àB������(vTr���6���怂��&�;�Ѷv�&Q�q̼���C�{�J������`�0�2B؂:��%��*]|�Gܥ��O'�_��P�r?�uOw'.,Z_.�9~f�-�M=�;�'��&�a|�ͿA,���y������ǐ\)�U���Ԏ�A2:�jD���.�XO�̼\A�5N��OG�2��uLԹ+���iy]�õ�ic�4t�h6׾����x內t���L���mK�9����>�sN�8U�:.�9���|�Fj���5�AD�X��D�q�/y��p�� 3F#k5���dٶ\I�)E����iI��Z�B̚+]��({�$�F
� �(p3�;�F��3P��9�w�L������*�HWL$��������Eq���O~�ޚ�ɒ8C��l�	痎,������^3�x�p�`�iSs�np'P)�'�6����5��js�큙�sDr\7�E����ǎ�K����X�k��c9��1E��jl�4���y��S	[Y?��x�/�AVW!0�Ӆ]�űx��O�ī#�2+�S��']�S����>�ݍ.��V����J#r{���s .�����ĨW6�p�D��WM�,�����El['����Q�:�m�ge��i�]��tǯ��b��/�Dc.�P<Sɍ��u~�;������8��>��&����Q��]<���������8HW̷]P�SGyjXJ���\X�����ash`ē����f�t��h�~��fK��-͝[�{�]W6UD�:�Dh�s���%�" Ɂy�� ��(�W���w����~�PhLb� )k�i�q	��V�7��#��\���ϝ���<�����{��-�>´J�!�NB���f�o��Zǵ����z�	+w����`� Z���XC/Aw��jDT���+�b�U{�g�t���]V���x/�]`-}��@����v=�߀�ț�)����D��pr���2��[�y/�LV2�I���w�3��}l�؜m�g7��"%��<I%KBs1T��]�ښӦ�]����S��!V�c��9j�	���և���L�)�~�:��:���l ��9�=�����{�Մ��*�y���}�
_$��V�OQ��0A�CŜ�v��-�C�z+��l$�\���L�zT�Jz�g��1��R͗�\/���%�^��K
8@*�V�ZI�̷k*�	}Qz"�u��Ó2.�OMWz�4D[��Z/����H9�ƠE�D���մ��k ��
�d�󈄜�ὁ��C�·��T� f�s���f�+���D��V�L�xh@N:��Kǚ,��F�p�M����,R�N�����H	�e�vP��RMJ: ���V�o웝"�T΀�)�Z���
"��[�bEf[X�/�R����[E%�����uf3���Ym�Q�w�w�,���@G���+:nc_��/�&c��?l���8�o}��H �q�y~�gY�sf���n)uK�����q|��P�z��ǟ��B�Z�r�b�O�t��ud�_�ГsFWc�*��Ӈ��0�����7Ue�;^<P�5G?`7�4�L]�BS���b��&�݅u�b&�>�,!>��=����,�������
��y��u�|�ε� S
π���xS��4��x���(q�����	�l~o�
�X��@ym'
`I_��MC�r��5<ॺ;��}:�v��Y��|/WWv�9�x矎�@�f�In�٭g@�6�������	B�tK6굀&Q[���u���:j	C�(��"�]�Xu�|
�g���m��򓧹�ܵDd�"�Y�g��%�C�լ��L�D���T[�'yrp��3��IkW��c����%ϰ˟���)'�S��}��Y +���SEj,c[�zjv����W�x�b�G�%v�U�ϲ w��?�en�1���XT<�$&&]�O ��C�2��~8��笹�ӸU��s`ܵ�Yo�Ͳz'���/�G�$�'Ŗ��J슏�G�87Lo�����m�o}�˽X
[�$(:��ݏ�◬�)맊�b��r�zZ�П��*��SH�l�g�*�sڸ���̫��(a%(�
~�m��6����<͒�nSnVu�+�*�DA�N�{�6�oh3��Ү〽(��ǂ@S�
A�1Y��
��ʹH��x�> s0�NA�U_PN�M�gL#����p7f����nM?%v`ٷ�k����b]O����*���v6�9�S��1:�/���O6sx��]���r�=A�`�N���NM8���1�/b��oՠ WIjn�/���E���������j�0�
Q�D��0���2�Y+��>o�`4�|c�����Y��IX4f�U7��/��@i,�/�N���/�77�c�����Tҧ{�Nn���i�B^4@��0CD4Ƴ�:���:�[˗C-�y������Į�^�T��Mu0��r����'˲�P�r���HLۨ]�-�������sar@��{�T%�,�b`I�L�.�$�Mx�b���@TP:�L̳��z�q��7��Z���j��3
]�~��+�w`�o���.a�|��JP�R�1��P<>'B��L�!#@�Ĳ�
ߚ乛n�+=�3�H]���e�ik&Ď/AL����`���Σ7���ė�	�z�&Y���%2�O45��X�F:cm�!	-�8j`{�wG1�W���ı�֘���\�e Hݡ�E1X-%�Že?�Ff9���A��?��7`lN�,���!D��Av��xd�E<]n�~p�@C�7���rլ3�K]�+��<!".����}#H^�� c�޷��o�c夻ğs�O��`��� OH�7(F�``〙%n�w���B��@����͹�^�V�<2�1�ɕ�R�-"��M�&1]��.tr�B��ڿ��Az��)��c�QAxG!��R4E���6;����v3�!3��o�?�"Q���EB�bm��٭44�c4I4��2�1�C��N&������7;r_>���K�/0���1��ܤe��f~> .��yq4�}��3nn(�8p�r�������sz�{0���˨���1]`UF�fYJ�q�{�x+
倁ƩׯY���L��!.xZ�m�f��ఓ |�{�����s��[.a#��A���	�@$HB#��O�1\u����`��}�U�1����RZ�����T�u�D�4��fc��h@ގH���v�r��ۻ0�Ŋ�ٮ����	��4�_K����g�_F1��_�tܮZ�y����y2�F4�H�*��K<����ێռ�D:H/�\r��o+g*�nT���ǫY��,��L:p`�n!7 ���\u�� I�mn̥�`c��B�KƓם5�̃Ǐ.���(�m�W�|�qѸ�e޼��RVW�lL����c�*0f������`�~YL�0�.r��L(�p�,*�<��(w��������%Z���gXP��n�}�q�hBj/��	P��Bz�g�$M�
W�*7�Kl�����laJ�N�C[L��;X�ꬂCq��bv��8<�W�vOo/mqќ:4�}���jL���:�q6�5�=Q�e�b`x�
��Ib=œ�jaVr	Z�[�I�tɠ�nz#Y��t��H0����%9I�,���8Ӷ$�n5����8����@`�z�		�|���`�W� u�&&UsMj��B]��P�F�~Q�3r��#���Ըg$oo�(`W��6fXlxVHYEB    fa00    1880�V��BF�M�\+9���8sT�����_+.5�e��Y�C��Z�F��qL*���u�ĵB}T��2� `���/<���36�R�?<ܩ4Иvz�I��6�=�3H-�z�V�Ed�[.ĈG����n2�\P*j�}�6Q�xS�%15���#���0<2���i]�Jƒ~8����2�T�G�R�\�r�Rh�T��NB#����~xs;�%6A�Jax��#�T��vr���SbKo�V��<g2�J�@���O<�m�b��0��Z~v��!�Ax6����*�h�z��ʆd��j��'�-PP��-$G�����#I�B����#yǀ�� k_D�MŬ��\���;���&��A��2��KS�p��)�f��,��W���_��U���G{dA�,n�]�"�M��Ug��i��7Д8bc����}����R�d<�rv���l1;�g�\!��*%L�`�A���){6g���=��x0�^эMu��]�֑N۴��ҟ#L��G��LŚc}/D����-1�����n�o֨:����X�����=���� ��V�63�RlS}�@C�^�vC���(Bw����}K�(��Q��y�=�&H���5�s	����
q��������ό��(
��	�h��K�V|W #����_&7�,\}y,�V�.�i��F�$�5ʨ�}�G�c:���|�&Z,36	V(f�;�ʺz�����G���R�+y�`~mx�_���C�L#o؁zc�.�Q#H��z���L���y1R��?Q����qt��!Moy�P ~Jޥ���b� ׬XO����FRm���O:�#۶2��o�%(��JыK�=#�y\�D�iA���R��5%�mO�ٟ&�&���y�a	|$c(�s�_׫U�C����[Z���8ט@䭭F�E4���M����.y�!%-T�6��x���Ze��x*�??9�c��Wkh�':w��s-6�{���IW5�_�{��]w��6�"X�������*�����D����a��Zx�`�Z��r/��V�%M�z�����C���1���� �K� ��Xt���Lu��*��A��[��)����35Z��V��Z(1=���Z�P�GC@���%�hP�����!v8�Z�O� Jma���:����;�뚱>�i���o4\	D8�C�0B�Zl�Ĉ����ڗӉ�R��нͶ�Ǹ����]���Զ�ŗf'[����� gv��ɧ�4�����s`���U�u�C��Lㆉ=˱:�Y�5�:vã����UI�?G�@.~{/�mS&�oE����15T�T�Tu�g	vƺ�$�~M�ſPkn�����{�5��Է�]�a��ڳ�*�����~�6@ɳ�Da������R!�MYU��:%�W��'jh������l��j��������|��H��@��|�o`�~�/�����Έ��_[���6ٖ"E��-��\�0�D@��)�Ǳ��!�۲`c����s>�/H�O��G���t�͔e�6��>�H:���-����,lX�������e���Fc���{;��g��1+�>�m��Z��&�t�ުy�Z�9r��71�;')�=�`����V��Ҷ�H�>���y���N��4�Ѷ�]��d���/�F�SOfKx�s�'TFe�Sl0$�D	R]��gn�OG+'+]���e\��L视m��$Vt*�a�[�V0�}�Tŀ�U�͓�̓xu����`�����V�1kD�K(�?��Ry[�~�y�����{m��y�~���e�N�_؊ӡN�1dz�;�J�ܫW�,��m��W�>~�oj�c��'?#,������&��ݱ&מ�D���i�@��OK�D�:==M+�?�CH�V/ᑾL��KS�K�h]Nɧ����?#�ҵr��*�7���1�Ϩllw���OA�v�����s�����Pqq�o��F0���PJ��}3Ɂ��Jd"�=1*W9��	�G_���j�/N���n��G�G��&�Pԛ1���6�w����mf)K~��#��`zW��؋��;G��Z;R�O�t32W�j���M�B4�lk�����PI/�ǺV���E�H7�|��	ُ@ʩ��d���M͝"�������D2($���S�9����m��'���qQ�*����m�m�e?�>�X��pMvB�����ʈ�*�`�]��L%p�����BLW�Ò��Ϥ��b5�(6�Q ���WB7���U����*������#�5�p��L %��+MwN�]15^qE`������wy�蟒��7��JX�s�*(�4�GD��-�G,j����N^;�D��+~����6�!<<EN�~R�u_4�+��ܸ��v-�ɍ7s�tŹ�����ɔ��ǿO�d�hM��x�)�#�(�O�桚!���7�9��͔:ˁ����C�� (���IY�$���`p�UU��_>�KG���i�L\W��@�*�<�'+�����g�hd��-���HH����̸�{��-讶Q�aS��Љ��q�w,:�6.����ࣣz��d��T���]gE�9!�|��5=���l�CL+)xدEI+�)�<��[K�3�tO�m	a����x�,��Z��w��M��ƈ�G!x�hsF(��`��S�&ޘ�\�R�l�o�����3g��M�aɻ_��XTd�;pD�ڐ� �	��f��;��M�	�}��G)���^`E���z��);#�Q�����ăP�)j'jJ�t�h��k����Y L;.��Н�����i_�Q@��?"5�5��ߘ������Uh�TC@�1�S��Q�Y��D@D�]�i`EG	G���8P�uZ�̓��DʭK�믂ƃ*K���m��YS����ؠ�L�>XZg"{KGYi������Ӧ�7y���\������[�E����������_��&)aeQ��V��g�\s���ÿ�����u1*z�_j�g"wP��5���g�H�l�Tx��E>��.�"��5Os��;$z�ˤ��VL`�l��}��[vt:�F�&��t^t���)*k'|���c��&%{�����vw_��َhX��圙ݍI�؏��H.��L��$��Ui4^���7<a�j3�#=�n6�<����;E��De�1��JS`nʊ�T\u� �q��G:�3p�
7:�QɰB�VAp��ę�M>�M@՗i�YC�aku�G���d����sƛ�����t̬�AX��f�s�̆a��!Vwd[������A�R�* i�<>S�JDS52�wI�洌%U���l����O���`���X�w|Dc��xd�hp8N�������
�=g#�T���>"����l���4{$W���z!��i�]��B�g����w�N�Ӟ�����<c}����C�jz7�Vtp�{��jiy7$��U���-��B_,��=��O��W}Oi9ۋ�]�f�ϡ'��R�%����$�k�R
�P=���j��G6Z+��M����䩄y�u>��Tu��ە]K�@ؼE�U�!Pu�f��	@-����^ơ"6�1�_q�����P
��v�y�7D�0�D�^b:+�~���ML7D��7� ��_��ʭUʷ�I>�e��/�)���g��/�[�k�/�[��#���̫�,���f߭7�</��%7���d͌ו��QM��:B�٭�'M�ޠ=�6��n��	*Y"�C�V:�@}�mqʨŇ!ާ��:�o�Z#�6��.Xܪ�_P0�v/���H��w�"Q����>��yۘƨ�Ċf�}>�.>֜<�	%�[����"'8)�����Rc�q����b�'ll�kO�tB�J�'e�}r��_�M�luo|��?�A�(&z@+�r������`��c��Y�ZERK*'l 똸@�^
J|h�ٺ��;Q�E�+���0���OV�-�U�\��l ����1�1�H�F�
�{�a+d�Z���mv���@���o�A؞In+{��R�/����+�4&7�m�>N"�+%N��8�A'f{�����CB�r���f�L.�Pڜ�=�+�����{��rD�#dי{�tL��Re��|�wU�T�֯���&5�RC�����gRۺY�����1"��u�CKn�8S���+�?���/�+�j&q���L�)�Fػj!�/��xP�	pr�19��:0Y�dCL�!� &��Pm������#�0��!Aoݹ��f ��7�z#�^r²���O-�#�YX�9߿��ּ:���R�׼����D�N��L��1��!��x]^%�R0G�$C��u�xx�f&��^�[xxr���M4Wt7�7����C&̆<��֠�T
e^�a��_r��Sǧ���K4&��.��*��sg�X��8}�O2f��.����F,�P������؃�>��oZ�TЀ^�R� �]���'��
OV"�[�^�yz���(�0[(x��R���1�B(�1pk�����������_�yS��tQS �z#J��﫮�O��$�©���:6)��~��G����M;K�����F���X����d�}�"����T`���*�Z �x�kv�ܡ����1o���1:���ds�>��1�tyy���^Kr�� .��1U�;����V���>p0��{��LØ�=)�d���a*v�#��j~p(���S!��J���G\��)s%�g�L�$�Ǵ&9���vb��x�G� �DǞ�5��7H;O�_�>���m��>��XHY.�&y��#͢�"���0�G�^Cw��b��'V�������P�Ũ,7H�s���M(�h�-��������2���D`��y��
�p���m�mj���氜ݡ>�xe"�UE�5�o,��0�wU���W��M�IMu94ݹ��*�T���y����P@l�d8q�.�4#J�T�W�F{\�5������I�XT@��ӧA�h_��O
!0h��Ͷݶ�������~�:g����t���h���J�B_�g�?/�|��"�I�V�q�9�߁�'��m���� �%G{`���uf�V[�������0ͬWaC��슜LWo�	倎�0\����V����%�U}R*;�k�����5� ©h༡N���!X�bv7�.���1�&�h��G�&��<�r 4}���}.���tf%�mo4���˺��̝	��Q�o�_�m����{�Q�D.�<�m�l%�^��+T��'g�HQ�?*�܆k�\�z�Vډ�I����B�}6���ǒ&���L���O�k����|��u��TLV
�,�[��0	�4��7@��0�&bQ����oQn���k�m-�O�vd*���krA�w���Þ���6�/�"��M�?�4y�뙍����#Xl�e/��sS�����^P�5�-(�'N�K �B���[��ݭ�r�*��_a�}Wg��t�/hXoE����z�Y��f��l�b[��_�r���֊�&� 5���n/0U�D�l��u�E���|�*D�[�x�����Y�q�&J!:�j*Q�(Z���eN��U�G&ut
6���F�o�92��{&'ȟ���۠A�*ۓ�ey��j�n��b�7p^+D��T�s�c^�����P0J�e�{��Xv0e[�zVƃ�H���{ Ս�P�:�OC��	�d��$<���~;�?{�τڗ��ͻ�y�qx�;�5��y�Y��U�p�������x�zf�ֳ�	��(�7����l@_�e�ɪ��&��J3jR��ȼ[�����u<���P`A�F��e�n+-���殰 ֛�ب�EA��u7�|��2�$A�Qz�9,ˑ���K�=F��vRpB�V��-���定Pn��,�m�,;ls������ a������ZcR�{o�,gu��@Q9_[�Y#L�Ďݹ�w~�]@sS�� ������l>�7O4�&��Q��Z�'Mʶy"�2f�����V�@''��-�{����<W_�������zd^��o�o�_���������Tt�:8p����}����K-�p�k��z���{_F���/k��&#_b��K}�?w.svu(��P��+��_P;(m�U�����P��^�k<��x��$$�s�}*�x�T�}C���~�ʴ�4/��R�;���BiXlxVHYEB    fa00    1910��)龔�,`>R&�j�y��ga�	�1���b&ՋA���Qf�gy^�og��%��cf!俧}=�"���,"P��G����At$
OODa$�]Ȭ5���@�gy���.�eȁ��%�"j���Y�ʨ7�PC��QXuw��y�T�o���~�G�\v6�
�7?�p���bkt!�qm���0������o���<�NY ��M{���-h.�Ӑ�!���ȃ���\s�R��y��s0�v���6��\���D�\%nR�T��b�E�_i}�#���)�$3������Lm��]Y<�]2َ	��������GK׀���Ώ�~�l��x��+.�wV��������5�2���~�'<r���D�
+��Y/�NOtO�Jo�zp�*��Km��;��M�C�� ��l�̴���i
�^�i�2�͟�G�6*��C��3��c�����8���ͪ=t�`�߂_���m��8��sBf{���S�7�3��}�2���~�0�=�x�2`�K�8M�Xb�q��� J4������ե��"�aO =G���)��!��lK�6Ku�d��T�8#��$��0��"�챂��۽�ΗB�.�¨��YO��F|\;&"T����WTy��v����[����+\�.TU�n��((2�!��O��@�oy�4�y2��pP�=Q�քY�U���0��� ��00:���N7�7y�w�\����5� X[��8��w].ާZ�,��{�j]a�G[��M���b��$G}Cow&�������7o�b'��&�$�� �R���jZG8Z,�K�.�ݭk$jhu*m:� P�O �бu?E�_yS1|~��T���UF�p~_$�Ŀ�h�6%��
��AI����iBC���G���ZH.�cb���D@��J�,����B _`^ �j/b3%�);�q}hl�T��
�-�f�YnV��*��b�h����kΡ9����4��̹�r�{��j�N�eG"��e`%�rS��J�`N�yy)`Ec�W�����ɏ��hW���C���3!���o������2mV�d�7���5�H��V��ECA~81��h~�%��z־�/�kU�-�H�@�;��T�^&���M,�K�	��s&�^8_y����+v��ˠ@�̞x����
m���Г�'
�ɝv����c��цqb�[��a�pC]�Ho�6��vKv��j��O;$��Kb|X�7�q�cט�d;�y�rS���e��Rp��'F�Hz�Op�`��%��5S��\��̼�)`a�	���_�|��z,_�L7��3,�m�̷#9m}�8�Be�#9[�J>HB=���S��~�6\fP�v�&�C�Yc7�� ����G�B~5�iy�ܪ����A,�v�VIyX���ev��i��e(S3)�W�FD0�=� Y��#����?�B��;���d6��յx޲ff��<"B���W���!��vUp����q� N=�*"�6G��gi������p�����.�Z�K����bq�7�iZJ��5���![e�xo�D�u�l#�r1�Y�:�>D:���rI_�S	�DР5���ԇZ��(8eK������a�_hT�V�L���p�`�;�KZ$��/��ݴz{�ZX��:t�^(��/��j�7��wׁ�9^u��&PMK]Ç !��86���g9�X\,�h_�����ʶ��"DPAY>�盶4�������p�;���;�zn���-6�2#�t��Ѵr�u$!�;R��H��>�J�G\P�����Tn<C�c�&�^���r��K�H��i��y�3D�mC��EL�ʘ�c�_뻁,�+�K��c�M�ѩ�¶���y<��Jjҙ��o2Q�L�������ur�V���}�e�R:$v�M�W��ӔӕA���P��6jIjګ����Ws�X>*���!w/W���8�*�ؒ߃�L;o}�����{��ĸ2�.��H��5j����+r�~L�",C�)0#����R�rt�*�S��@�5��H�#v������|y�!Ռ���t:����wg�B��=�d�� �JuڍK�y~ٽ;v����&)��붆v���⚈i���X&�g�����TuwR�!;�iyM#��0 /g��(Q�_%~/`E����"���ܞOz!Dg	待(����Cj���W&������T��=7R�tˮwPW�n�4�[=0��&�/Ru3�=~��!{�'�No˜\�q-��:�t�A�����V�G��*B��� �Dj�����6��ۣ��f0��$s �[~��ږ�6�	�+&���s�߲d{��&��>�ə����J<gZ��Id4&D3��d���	AD9Bg�6�>��,�5����k/��>aa�ʱ�#������QY��Oo�4(K.�ȅ� ٕ7�*6J8O�~�o�����s��>M�4%~&��2�������	�s��g�zlКdN���AM�[��Q�&�Qc�m"��0�*k�mA�U�Rؚ -����*n��*e��y�߭r�J_����ޏ�������"J�����̉D��o?^b���)�e��$���C�b�Ӂ�$,�������Y�ryW�6&��+v�)�r�'e���D
�1�L������0Wx���U���+���\��UĒ��Gm�c�1�ԟjO�~H��xGt�ɮ�Y.L&w�X������|/7����.�HO��9�1�F�O�X���J(_��~��-�����EG�R�"5�Иj�V�An9�-&H�@+Uv���Z��t/��Æ�1>~k�Ě�����Oq�͘?�y8h���>�b��^�ʍ�ߕ��w?�>� �Ņ�Ұ/�&)��Vl]+���EE�T&����*�D�O��:��hy�2qU�W�ƙ���o~�?6���l�����F8�L�`~r �1?2}��c=����!,êO�PO|���?�0��~���W����rQ/S4�3�y
��(e:aWuj�x���K��>�n��� �u,���n��S�a����_�.mGեН��Gq�M�
3Jm����Gu�C4ځ�����6�\z����ߜZ��n��y�'��Z���ER&�2�4D*0r��5���In��b3Ǟ@�	�����s��N'��4���1#�=og1[��WYv�����h�#���Gl�����
H�̴>��&]��lwV{I��!g/�/�sԞ��x�){T&9����ݾ����U���H�� 5�H���{��g|Q/�r�Y�A�,��V��d	��X	ʷ�!e��=ۍP���� ����wo����3��.���L�`�~�H,��1A�iL�T�R�g��Fȴ�3M�|�Y�B�#0B�5NqSv�y�d`�¬���s���!�;Â���F����bQ�0��A�C�.�إ����78�{��@+|V���<��v�6<G��$hV��⍜ ����t7�����~��p�h��w�0�?-_J�B��Q�,Lw������q@NW�)�E�����!�S����/_z��D��@���Ԓ�bo�~���~��35P�v!�Ѳ�z�����#�j�ۊ��5�%��'i4�/�#$��LTp�Oy�i��iaSe��1� }�����~��5��.y�/���O���ed�ht�#��ig��u&">�oB���fҼnG��dS�g��G����}{R���QA�r�W�ZBrK�� }���U3ռщ���A�'p~��闕&5-���
�ta��4��W~ �v�	�K�XZYv�ᆵ)�=����)�+�C,9��1�va�q��e>��Z ��5�9��7w����ڗ��[ߝѰ �!$7m�`5����@��|0�Y[}'�s��:f!N??a��&g�j5L�*���v��"��l�F����ud��2�x�&��|ŷ��� ؉��?6NX�-�ON�{2���dW�լ ��-��˃����
��m%�?)Z9T�t��;�DJn��X���Q˄�C�QDk�A7�{!`T��4�@�o;�j��6�C>^�v'��k���>d�!|�̀kC-��ug���l�$�w����v�.4�Uu��-1ޫ��~�>�S�����	����]���7W�_��.��i�^&F�����F<Q�Y;.�_��d�����*��'ZA�	���b�n�L���evRSq�랛�2AX�
) oG�������~��Y_ ����e�иw�f[r�2���Y	��G�Z��n�kzT��uZQ����ŉ�g܋~��i�/{O" ��Os�U���Dg��-n�m�ҽ�?���vWm9NAAs��~<�^l�qU, �|�[|�g'��5H��Ր���4��sNWPk}��`w���3��+�����JFgy��.�	��s�!9�o:>�> ����Py��ۙ�+�������2z��Z��~;Pz����2Y��
�����y�g����jړ�ݯq�@wu������&<�������v;X�e�$���0^�N�S�t����I8�^0�:��w�h=о��*��Ϻ'�9�ZI�~����b�y-=��(�LJ�UNao�^fRHk�J>`���?[��uU��v^Nζ!h=��ŷ�Ꙫ~72�ݸ19hڏl��H*37h	&�W�UO$Z�E~��K�};R��`���޾��H�-r5oM0�" s\k��~�]g����*UTD���_������E�p�R�R�~֣�������x�ev���ɻv_)��hW�Y�g���G״ۻvi�¶H컕��Ւ+յ���>39�C7�^�+�˺�z�	ȁ�0D�'#�5W]I���X�垣��hS�v����I�M��Rm]��2ʄ~���ql���խ��e�{�Qv�����$�3��k{����4��j<�E���K�T�0�N����2i��\1zaM߶)Q���&,���L-�<@����v+�����IK4�q� e�l����K����*����X�e1^-����N(Oـ�(�7�8���,�2�\� 
S����W��d+1H�n��=�س-[��7n�x\�S}v7���/����~1�T���&\p��p��m�b��Y|�1�oZn ��o�i^O�=��8	����	b��8��oK��=U�۠V�4pT�Q{�P�K�G�^u�ǫ�������^�'݈��|���-�)�A��x(���=������ǹt~���~D����g����#$�:ۅ�G;�s��e8d��57ȶ�(T���S6��h�,��:�|"Qj�����ui�`��ҼZ�%8���&;}���,$��fn�ܴy��~��h(8*B$�#?L=i�m:�J��eKɩ�`����P��`�����o3X�nЖ��?mJ�^1��9�n��S6�k�����@akJW�t9a��`i��8�@���v�ؕ�UZ5�X��
dF�8�oR�`� �޼?N���x��Êk�;#p#.e5J���N�Qa�ځ��`J��9�4"ZJ����H<u~$z��p�?W��&8B�aC�1�$ܠsfűp���h ��:6�E����o�d`V�V�pS�1gȦI�teMo��/;��IL�;w��o)7��]0,��Q]�l���	d(���=�z{�A+�A�"���q��WIe���TƆ��;C����e��\����w���`n3Y���w�0�t�*%��N5�/-S�OC�4���+yBL�{�s���Hs����)����?����P���k�IG�ߣ�3�e���f2@}��?4�Xm�X�#pE��Nf�Ldf+Y�u��;�bQ���vY�ʐ(k5����BSK��'�z`ǵ�1���J��¬�`�T�w��$~�.��Τ�g�AT���9�T*����z�aZ�p�����U�+j���f�3Hȗ�S
�r�fkiO�։��;����Z_W�i�}���c�R���{PD�I��D��,�A]�ͳ=�]e�Ԃ�G�Ϡ)O�\�RB���/Sډ���g�����"���I����Nu����n�I�o�+7/� V$����1c,]�hf����X���~���׺mQ�.�����*5]���'Du���g��D�����w��R׮�4�/6k���2OQÎ^2D����_`��}��P��j��
U*��fޓ|��NEch�#X����K2��_�F����f��*o�6�_��!���z���,����n������ d�CO��]���F]�B��yR�}z�p�/���Wa���G�,�|���;�[c���zz�*��Di��@�ä1���k��XlxVHYEB    fa00    10e0� t]���,dM����QG!S�e]k�,C��O1l`M��Qg�p��?h&�@*�[PT��2��y�{�o�{��AM�q2=
��VVΎ��=~�Y}N� BU�+�$�1�}w�K�k����d�*a�=E"'y�rTL�W�Tw�������d-/lW2-����.!C�`�a���)n�Q��B���e�pv�5�_[u�wS��>��d>��g��'�11��z�kՀl-<�8Ҥ�Ȗ�j?�D�Sx9�+�:��AP"m��0�}����y�>h�i�α���;څS�dN?V�$-W(\9}�5�{	�\��7*$��
a�<��N?[]d�*��Y�[7�򐡜}y���c�y\�Ɉ��>r�X�;�:�Be;+x׳�5��7D��VY������6<��]����1՘C��72���:Ho����l�ƞ@���6@2���w_1��=��'�O����!pN����*It4�k�GϷ!�Z���J#�T�J���%bT���[�Hg#�I�=ރ,���C^�r���QG5���+&&�K?F�j�(\OEo`�BÌׯIyqEپM+�b�
��2H,Y��3���:���h�+���>b�!�-?9�u�[$�9�D�P��l=��+�*�6/-�0�yH������wQ:�w�������s9����_�`AZ�>!I�[؜$[�qNq���w!�&ǧ$-f���[fN5
�	hz�x�5�s]_c�M:aі�p�a���V���Y˂��U�Y�M��C�zs��Q���&��w�����	v�G��{�X�@Q;��cS0Y���MP]�s�Y�>= �7��S�5��]��v�2��fLy���Wˍ��ڂ�o�*��҂� ���يL-q��l>� �����Y��[8������1ڌ�����:+�6`<;���vC%�a.>��B[\b�K�������n��/9�˿��m�$x�i�OFӢ��@�Ϳ��%d'�Q�U�z���1bG}��/��J�1{%��!��ՙx�H U�+�0�4ނUA���W�^��]��p���Wo��g��"U|-��m9����f�t���^� E��KɊA׷�ho_�mObu��4ס�Ts��za�
y�Q�M�Ћ*�֥n�0�NA;lj��^���q���Q�WovBwޮ��zkFY�j�\��=)���_�fٗ\�k�t,��-���$/igTZM��mQޢM�g���?`a}���oY����xK�F=��@��S����D�t��F�F�zH1�H�)���>��&��$�T�XQ!Djm�Jd,��K�DVm4(|����s��<{["��W�;����n5 u���Q̹���_�4���M�k}�8�ˌ����ΠҞ�ݡ5���M��렙��'�n�����{şq�3i�ݐ�X��bJwlR=�$yd��?� r����t ��ȓӯ�i�������%�"G^�*���ݷ��k�qnt��ٔ����}�UY��l���W%2��)�����&r�O37�``p��&�B֌���^��4�b>��%��][�1MA��h ��=�oU���YƝqp�)�RK������g?I����yB�hwL*�S{(�O
@�e����k����%�:��xRԠk��۰`�^��r�9Kg�)��s���S7��9mP��Ae2���tSA�IYŹ�������Z�0P!$2A�7p�<x')���̶W�˖�2�����8��L��q��{�V?Ma㬿�>�r_<����b{Y�/��T�M��V$T4l��E5*(%�d[z=��`(c��;x��h���A0Z�?h�0�ȯk�\���Tq�{������*��������3r�9�C�)�hvp�`�%:U��@� ����c��x�b\��M��a�$���}�C=�(kP�����tD<�UBΌu�v˶������ڪ ՝zWd����]C�v��.���+s9����� 7킘��� W;�״:�}���33 �t��C���	�9�g�_�ΒjboH����I?�;@f(�x�p�V�6Nt�'�U���������*K#�⭟2�}"���<�ؙɟ��H�t�r��(�x�t����>`,���m{�Ib�ݤ�����Q������l�P�(��`��{[��\׳F���(cF�)U��v�6�ko�%cͳ��
��_Ϸ�j�j҂��`V�6��0~��"XKB�?�vS���Mus�%"���b��.4lב{H&"��Ci�4!6��\���gr�E�zG�����-X�50����}}��A7l��0�T�G'{�Z���`b� ��Wie�}��Sm�.�TG��d�"M�y).M5��C6���e�o�Ml3�������!	p_i��H��7��CȦiB��Tt/�.{τ���"�����t`/*-���O1�*�x���y<ڎ��N���D"�5|����_.�r�NwZ���Dq��JqX�U�Ad�j���ɸ��]F�ڞz˜-�sN�]�	�)qz��=V'�n<�R�����������v;N��=xH��)�}��kJ�����lf�PW9�"�����Y�6Bza`Z���Ã1���T���Ȕ�F����������tM �V�9��b�������_9��d�3�L��8Im�͋�'d�b��⮸�����( ��*!��X�{"�Y�eI��z%*<��������;�.BЋ2�d�"��t�$�Z�6Z�SNBn�u���I:�7�g�RwR���R�ԫ��bQ��VCĹ�t�l�����8��&ق>}�g���E��ˠ�O�X�����nEi2����4"�|߰�a��H�I!�-����7Ju/�.�ޯ����IPjʖ�n&��(����D�/~�K�M�dD��j�O���w�j������|��J%x�Z�f�ZJ,r�#B^+t����l(��R��Q]����\ą}��-�Z"4Y������{Kv�j5�Z�-��}�=�J�����������W�y�KAFxG�mnv6����c���Snf��h^I҈��7C��9�}=g>�����
����P?C��H%��@{N2G%e�Y�ay>���?F��|J��"M�,�d�d/��`?�7EZ+r�Y�����c��̋�O`��h�i+�LH`����uK�N0�A��Vls��0d�7;�-�(�X��!�c��{[<O��)ĺ���_&Þ��ʇd欲O�;��_��ybq�b��e�,{�����Ye���_v�;i�����<q���iK��<�� ��d���C�:���®��MHE[�Il�(f�	����(����1��ƾ5g
Rjnj�4�������91���<҈%Ӊ�iZ;v�.�7��䷚O��8�}U�`�ʔ��I��R�H�3*h8��(_��X{�n��O]Z���8���p<L������荰�n`�h7E
�<�%G���0�'���1۶�Eه�b��t$
ط^==�N�)tn�c.����4+#�`�)�����'��t�Ȗ������U[��R*7�,G{��6I�L�q 7-�� �x���L>�+}���F�{��]�OzBk�˛�ȑ�)���8�u(d1�}�ep1��3�Á_��#�_�:��j	?���k3
�fC9�:g9p�N�H�h��Sz�N<��ڨmB�ӄ�<�(�g��3{����~����3�����>�`�rG��+'��>[�-����z��1�ͷ�zKtbNoT��[Tb8��¾ؤ_����(NPn?�f�Hs#�C�z!�6��=�'���4� \B�1�|/�bE�p�j��	���͛�nq`���zt���$&22�T`�>Lt�W�!��P�F7Nf��nŧK�Uk�����A���!_� ��ˏE���2� �vDS�s�u��h�^���J���j@x�3�r��]�	��]�:�z���)���S���Nٲ7�?��n<O�g����#P���O�wK����[���ML�5u���ׯ�m����_i�Q��3a�H��@�$�$2�E~��0~�k��!`���z RU���rm���x���%J5���g�D���{���
ǲ������-�mw9�k�{9֬�"��T�^�¯� ���=�R����s��8�G��\D�;L�p`M[P.���2�Ufd�S����T��|��kӲ�! z��@�o��F�K~��ci��-hXlxVHYEB    fa00    1860�z,�2B1&y����j����O��L\߈;9υ�u'-�W��te���W����79�쎓L��K5�|������r�j�PTvuԎ~��}�G�{:U��'<{�М՜���IƼ�"���\/`HQ&��Y�(���1�l�,KBS�C�n��l�c8� �fo��M3�uiǵ��6"�_�����_������'�[>����<����X�8��
FF)0&_7���Z�R�f���' �����VW�v�]���߾�a���%����xv��D����U��P����m �������a�.[�1K݀�ՐT����Tt�߹79���3��X�lַ�p�b��(�N����Ljws��5���f�|�/#�nyو�;`��+�I��]��C[WH;���gP�e0$I�p�j$N�L����!�H=��� "F�N�ss������@�q׺���UU��.�,�����QoH�/�w��)c� @E߅�-��VH�w=�����{���U;����K�D��a�"�g�k����Ұ�	HM��H?n�g��k��BhE�	�xl�sKK�qH�|�{K�_o�#7\�؀BzWJJf��E�}�z9z ���*�_�*�f��@���j1�BXi`��5G���g#�!�/H.�@�� \��G�a6��E�9��?Sh6��^hG�"�"%~��es�ͧG� Y���*&���V�ѥ���C�v�+�L��̦���%�@͕�RH:)�92 �>��&,�/�rO-�T��������vdf�1���G�kh��<�>������KV�+e�/o�-����M����Hl�� �V���M��G���P���3��6f�4����o*�� �w*�^�2�|�nȱ�j(h��k�9W��}>�	�\;�c���3�T�9{���hf�A�E�"���+D-k�~Y�/$��fh�G
a����x'�(�Z�m���6�T���[�.���2k��y��J����E<�;r@޾�˹�/ۉHi��P{6����#	������PDK^����&ܾ�W��x�	�ز��{�E��U+|\���Af]~���ldL�4,���2B��'gWI4'�`a��k��7_ԡ�쓪��'P�7H��{�*7,�8|�a��������:��矾�u�=��;+c �?
R k������]��Bu� a���$����2���'4��5�C߆�R
�oCP��2d��;���	�>TLC�/nA(�]���b�K�3H��a���1��BG+/����C��B"���ͅ��^L�����(�wӔ��š ������ Cn��3Fˊ`���²'LW�+%�k���J�ѨK�����@1�<yl\��}���dSX�d
<�x�P.��.H>��b/�q|�9]�W�|��ơ��/��X���7��E}���Tf������t�5-���k����
��Vf�<�k�0s�m�ؔ�%�؏ �k�@p�����~���.?��}
�H/��{��ch����I�U|'Ǳ2y�;�M�4��vg1�^��<����5k��aH;�"D�/��D��1P�ٞ�sB��Kx=z*���Z�p�!ُ �sF�_z�*�e���t��[�ԎF���ywH�j`�񬡷��k2�T��.�5転u3�K]���~��H����������zǆ:��6�O(Gi��O�[�j�5׎���<ȃ��#Y���.�4�mB�)�6ov��s��F_`���X�6:�'��Ug�5���.�m�?D���>�}�yn��~YVwX[髲-�/ �B�5�
cˤ�){=�x
�m�m	.��b;J��k��#6}��8Ӑ��OZ�YS9/tW�~s�O>~"�l�B^Sg���9�����Fݱ�1�؃+΂h�Tݮ_js	�����'dY�A��=�����=KWzj���(��f�*N�KYO����O �YJo�R�v>C����x@Si?+���f$����i�S����{��*!�H �S�E��E��K_OܓH0��W��c�Ԑ.�[>�OE����hi�H�ˢ�����o< '<�$-']qc���|TWt�c����2O�����U7���
d#�ӆJ��vJ�C��ϱ��f/|����-���$�4ZO|%.>)����L�E�T�	��"�ѡ=ыV�#��dL��4x<���y�����s+�ɮ���'39Z�$�8�f�F��,}.�B<�w^�<�|Պ����Sf��ߖ�A�j�*c�E�?Rq8��B4q�w���88�s0s�bk�m�}av��X�o�G0�]~+=6�=�B�������T��&/�v�[��Hi$�4)������l�ړ�x��<Ri���Q�F���l)�&Y]j�?��K�g5��s'u��[z�\�^���@B��֙~�הįVp8�3�E�}%�X��y���m�?�!b⮱"Q�:�M[�tg���:���H4ƣ���GIA1��A>htq�
��$������c&6[��;^��A[�#腓��9<���O���MJ�H �-�$)f���0m>B嚆�I"�O�f�qR�<g�5�"�P�#{��m�GcR<E�jxzӿ����
wr�7��l�B[d�}Z�+��(��~!���GD���b�v�t��q �4�8���E[�
���^fL�lx�w��D�u��Ŝ\|�s��� S�6��i$a~
��,̠HA:��{P��jd����B'�XĔ�0`ZB�Ȋ��U1�qm6����	�=m$�k=S��g�AK�p��F����l7n/�ß�!�E��X�B���m.�ږ,�|��5
^H-m܍�Tŷ�kұ�m�`�X�<�K�{gy��s��a��ƈuz�����sy��Y���v�M�C��,?Dv>7'9��^��m�t���F��hz�P���z ץG 6ܔ�S��!�I��֊xLP"��������>��'�X�,��>i1G;7Y:>��;o���^,�\MM�k�o�l��g� ��G�������Wp�G���7��Q�9w�:2B��Ege��Qݞ�'ϲ�E����?����e�x��Q��N4�j#��"��ےH�3�Ac�����l��>9W�/�v}�?��"h�Zߤ.�*X�ׁ��b�{{5�1�ץ��H��*����Y��}D�/���GA�����f$�S�[4x�ac�bMR�})�4��e��
�)���ڈ��i
	���vM����<
Ϧ�m�7@��	%`Ʃ6�������f�5�:d�e'œr�఼�K
�ɔ)=fsF���;U��#8%M��b�A��6�bP8��3F�~5O/_������E���򶠷K9>X��74o'%��*"��T� $l�7C�{�O&�y,� �5�ބA %�����T�d�|6�-U�"���u&�5V����9�gK�M{����T""Y�zO{iDG��[+�G�~��ӢN;�o����M|Pz>�pH�� ��
m�4�/���2�ӿ̸�*R1���g�'�ʿlZ���e>&�yKx��9���bDq�t?�.��=�4��h�E� ��Ҝ4����J����p�Pk&��eَb"��/�_��չ5�{�њ>��uIq�n����KE%���_��x��$�+��ݧW���G��6u��IH�/H3Rj�̅������F���O��J}������4���H����ҒҤ1����f㋋/��ă����1�J���OlJ�N�;�pB�R��/F،R�Y�L��$�Z�� G��@��f7|�wY6w�՟W��γ"Z��Eʦ7�e�&��4��I�M�؆��;�^���	Q2E�Zs��R�J��iy�Ȩ|���m�4wYJ9�2h��<�z{ٿy]Bd����/c7�k����^��`��5&��"4��k�cS֏Z�|q�V�Խ�Ȟ�Z�f��]�\dL�J.��=�ʬ]�K)y�[�.���#B�
g�E�����zj��F'b��K}_v����Ds�dѯZTمpӲ�&dP��_ĩ��U�x"q�'�����^�5���7+W�}u��)�L��#P	#�^�k�_\*�!�Qtx��;����W��
[D�!\��+vxqp�E$����⁷x\� ��s?\�%�������K�!]����r-5
�^t�ѣ��^�J[J�8F
G���?����%X�oT��]۫�`1'ɤ�#�nj{!1�VUM�D�{a��qc�>�ظq�`�ra���iwe`b���+C�
 ��N{�x�=��Rj4�n�6�m���/��L��jb�CD�0|���?��t�U�3��1�N��4����<���9�B�ių����	+�aL�.~�	��g���c���GV��Y���(�>2XI'��#�Vu[�;�D]s���2.�R�@>G�2z�f�Eg�ߡ������9W¤t�;B��<ǝ�[��Θ,��6�cvnK��qJ�� ���FG�ӭQ����dM��&�,_E>*�;�i�94�#����Wݴ���{�5]l��QW���P�����R����V�!yC7�$�S����R��FMb��=��ONǚ�>׆�y�Fk�dn�>�m&�COH�3D�H�b#!z��r~���jXȗfVO��r̩�^�0����r^����3:A�d��nC�!�(l�)ڋ�Z8<�Kb�n�Ι�+��=��xۄ�Ve84�}�3��Q�X�Pu}zO; '�O5�"��{W|�N�	�U�>OI�����a>���_ڌ�~�D3�\�$!RSN-���[��^�P�I`�����X�o�n��{�%G�K)o�X��Y.Z�z+8�,�v�QV�3���2�~RRiU���`؅�}�4���`P4Ꟛ��K�V-C���z�\�/��ѻ8�O�{Cre��y�L�q�A�F�5z�:�&b�#s�@��C�/�7���3�\S���g�Nj���=����$���n��N���Yk�n>�j�?[`���3�^uZ.�W5�%/��� ��ӳ0y�|�;Zّ�s�.����첣	��=H��+�w��]j��Y/p����V�X��3��;��.�+T�$qX��Dr^6^�i72�H�$�ܺL������z���Gd�lp���2��
2���w���{�}0�1�PY�1��ڣ-��"��B�
�z.�W-�(k<�@�w�yȆ��+���Ti<��N4�`b�)�V�@��0_)q�9v���J��J㸗��r�֬
�/ר|7i�uXܔ�NF���[�ҫ>�0+yo��ޑ.�0z \]�=H���@O}���ǣfǀ��I��k:ÙԶ;H�xp.�% ��Ka�=�uVZB�C	n�%�xx(qo��4��-I)=�>�#��f<�s�WT1�G�&C�ƿ$�͍�DO���Y�YS���o��G��!�v�B���s�{-�=��GV��E�*x'�;�ӵ���.J������r�����xCժ����{�[�����	x7�yed}��ex�r�(�aP�. iBѿ�` ��4����a6��-�����Ж�*����>���#�=HX!��-5��5C���6�s��kpFR-j��ilIf�G�T��a	��cĽ��O�x�Bp�EzDs�-���M�� ��@򦴄��7o;�� 0�=����x����%W�øb5!�=��(dj��:	ɯ;�Y�=�8�'p�f�8�^ٺ�9�C�r���ǬpfvV'^��d��)4v=s;����н��%=K�W�8��Zf�N#oW�f
c7�d�v����*E�V`2�kF#�;��wk��!&#�eK4��I�O�g������@F{U�j���"�4����Epji!����,T�޷)���,v����VϤ�G49ȭ�i���L�̓�1�������
�9�v���Pز���²*��Xɪ�ϘQ�λH$�������X��|���#Nh�OTIy�=����b�����=�:�(��i�)8O���U01l��s];T�S��sh����p�*���Gȩ��ɰ
�E	����y}Ȝ�D\; &�D��t�ʙ��,��N�z��hđ�`�u��U~.��X"Z]x�c���L r����9��5{�bP��;G�h�d6�%��vts=��+f�� �~��+Q?#���&1�:p+c�n{��>�c���I�:�9>�����XlxVHYEB    fa00    1720�uˡ!-p��՝n3�f�yn�k/���oC9�ܩ��X�z�cY3͎�����r�O�ڤ�{s�:���SY��ZnQ��.z�8Y[hh9 <���+tT�jg}�S�Do�,�^~���*�Լ
z]��١N6�E%V�d��t�o}@̍��ZNߴ�f�:IJ~��=��A��r���]�$ӴTWp��%'=a���Ejn�v�(1V�/�wg�'#�4E��s���:B��
�"2g�|�EN�F����@c�u��� ~ �� 
T�oЏGs�Hb�׸�v�eX:TJ��7�L�,�?0;,���=��SP('45��`3����+a$��ܗ����[F�u���~���4�nV[s!++�Ԍ���������D�;�d*&�J?�M�r_8_]��F��@�������`��#�Y�Ԡ����)��dcIc�Y��VNȓ]!w
���^_Q�_ρ�/� 7@(�d!��*5�Waf�e?��S!K^X�(6}�OCI�O���Uk��&(���C�4)u�ڛ���N�o
		�z�7Ba��J���'?h����.�S�j���]�<�M��H��4��axNt")Z���V��A�Fe���1�?�F�Y�2J\�������@
��;֯��) sud/l����/�~����ώ���DG&�f�4NM-�lN�D5�7WB>}z�P���
	V9h2�6?����oe��k@ �v`�q 7����8�)�y^\���]`j� ��N*����?7��o��AQe�K�H>�Of�C&��l$6�ZJ�Rׂg�e2ٯ�Z� 	x�nMӮKm�A$	�N�qk�u�(�SCl�E����`�$¹}��CMOjԹc�H�V�O���C"��뇝�-a��P1Q���)������R!�nJgx%�q��*@+`lC-{�?��Z؍��ӭ����{r��vG%��̕(-׬}��5f6��E�kb�����j�F5͇�8D]�1�T;ó@�^��w��b�)�)�_� �����R�BI�[�E)e����U8M�����+~F�UN�[( ��R��a�s����S�@N2��@Q����{L�n��I�o\d�����B�1�����!�@׿������#�߃;�.u��<BB2 E#��BT��$� �������X���\Ƣߍ����:��՜����
���8c3XrwA�?��'�;��1�5��V�H�[�+dw�.*X�DXD	A��z� �����������U��� !�o�Of_*yŵNq�<N�Ә�	����S�Pu��c,&���)Y��%�4v:�1U	�qu&��2;����C,
�k�8ڀ�.�C������� -� �ᯩ��=�����������^�3�Ն�Ɏ�����gS1'/���{������c�־���)��VWPR�E���m/?��X3����?@rsDL���Է��%��w�ETbpI����^�K�YP�1�v1��2[�:�*�>T�(����s{<�<!��9[}�����^8�'��,]WҠ����hw0�]�~h�UaM|"vk�x1�!-k�z
ҋ�n�l����]�_�d�&p��n�������oM������⫳�x��oܗE)/�<� �K77���vqp*���c���0�G��d�	�~��:q����VW��2�]���x)�a��S�'V���KQ���̖�x����v�����_=�	[����Ex��6��*�Պ���� V�
�,�{�3+���l/SS�؉S��Y`�c�Y�	r?!����9e��6O��G���g2:tΓE [6̕À�4a�}ǧ2�n�g�����5����rO����g�1Y�-��
yr/Π����]V�Vm����l��"ʚ<K�k�	�O�JW�[^)�˃�K��b3tb�OE��4˻�[�d��K f��R�3�6���}6����Ҷ�� ;�TTK����D~DJ�:�'"=����ե/ï�	w�A
=��g�i��s�k
�g�?l��6_�B�[��:R�|:���i? �g;��%�p?X���[;�����E��"��(��_�t�@���h޽֬�b��}��� 5��B��ƩNMa��w��L&��U
�������.K��kp��Ⱥ�Y!���(c6��Q��e���j��"�3�x��u<�T�ԋI"�ڼ�������*k:�A���m>�4+���CC�8|1��[Eg�F7F�^��J��9�6a��6�O2!�	��	���濞�I�S��?�4���������eH�:h$��q/�Vh-�ۗ
���{U8�`���+���(܀h��{>�^�A�K/��>���
�;��`�����Ŷ��?�@�vЂ��j�_Lm�A�S3f���|gS�P�UA,�;�k!��N:�Z����/.[ [���-ȆP��;kDb�M8W��퉦��p��Y��[�c�*B	�*z�R����N$���,�����y�B=B�̡����D{/AE��B��&o"���� NH��К&sk��>9�8��%�w��3��%�G`Pf}9�������!�³Jh.�ȏ��n1D���QV��}�7�9\I6���
M�AQ�4��nɖ�L:�
[��~�^4'm���d'��H���y&T�<w�Mh��E��pH8�L��*��m��L�$:��Wy>Z+���h�~�X}�kaow|0S���	�	�=W~�h�q&(�˓nn�/�z����pΛX�K�φ��:,m��yL}c��V�s$H����ױ��J*3rt�I�;����C
5k�U[�Ȑ=3r�Z����'��t��nۧ�XN���_Ά��sv���	�~!;U�,$k;��`�e.����H�bf�B
���̶�"\P��{^��w��2�?,���0��HT<nCP�>~Z�����̼�%�o:\�'�(ғ�CU�����bH����(Q�P\��`��V�p�o&�����J�}g��)?)��B��8v$��`��E�ڿ��zlҕ�m�����k�WN���ֶ���L�n�{p��	�5��*r��81#��ߎ^��1����M��2�\��=�����bC�((���4<���ч����r	�*��gϪ~G�����__�_�v�/5�Da~3��F\zA�4^���H�Y�θ8��@�&ӫ� t9���M�diꕅ��"~1l��6͎�Pdw>������$�~�(��&��f0��~#|��+-��o�4�	)�6�|�������f;[�2��84w�"��	ͷOJ
&��~�l��|c�Ⱥp�u:[`�b,3=����R�;r�v��qE6�i��ٰ�',�8��x<g�6s�ɰ���7ay1��5�	�Fe��/q�T��3���<L���֎j�k������"���n�\�G���GD0K$(���G1��"X�5�8�zLm�(��a��7���o�>���1

w�|{�k=��<)AG�O��~/���HȒ��.��\���n5:�b-0���GA��;<�3��}o��!P� h2�)$�A�r�y4��l�gj�}����\�(�=ݵ�h����L�9�/+l���Zw"�V>�J>��x!oA@a%R�����x|�� ������Kv�Jqϭ�S�R���`����7D]v�^:N������t`@��Ao�o��](����!/�*��p�ׄKWC���'bA���C�����	�-s9)Y�o�5�.ٵ��K⇞	s(5L�T�Q^B�'P��Cw�'�l�kjO�c��j�Rm�#�J8Xxb(ع��+A��~ֱ���x[�o4�3�1��ȗ���kc�at��v*�	�0�8���M���
Ɠ�ҾWx��ͧ�Q�?��/՟�~b��e�����kp�ܟ���nT���CYz�:U%�`�l!oR����z�.�W�h�e�I�^���O���l��D���)��)G�c2��w2�גj��W�U��|m W�n��-�jT��)�����b�(�����	,��uQ6=�� �Q������KX��Z�@8)p��B��j���yi���i3��NE�ʇ�W�.re��w�����P�Ւ����7�0`}�+ȹ���x����wڨ�)sEF���Ki���Z���*픠:RR��]��{~c�2�1U[+Cv���z� ��Uӯ�C4���|馀�ta@2���_=��5IA���e� Ň��ń�����U��-�*"�������2�KtdD��9�йQ�Lz���=�R���QTǔ�SN�.���	J���ST(���W�-QG�Q�.���C$c8�`\{2hmE�<]p�T]y֭5JC��ey����aS���dX��Ms��T����TC�B2-3qs}�O�5��: {�x:�s��i�T�\�1�q�gr�5�����QX����Y4��)�����q�	3�H�-.����q~���e�ė!�ΦQR8}��H�T#ƌp.�D��{�k!��OB�d>���y�D"b~���s�:Es�Q��0ߔ�c�|Y�s���r�(?�)��	�/�Z�V8��u�)ny���z�*0�jn#�W@C�lO[]V���e��3��kt鉬����������X?�����E�����&�E��D���k�]� IR������ÁU5��y�i�
~�O������d�00���
��$�%��m�:{�
}��\"���|��%�T�����:�O�RѤJ�9�u�y_��ob��.�%[ nq=��X�9�4=��u�8@&����1��H��絗,��N�p�:��C���bB)B���D]�i(��+�bG��8�MBx��J�Μ� �<-�u���ٕ�g�>��p���d*��:9o���I�/�뫖���@y�.RλY�f���5P�?�)ݡ���Q�;AA`�����k-�P[ThI��������\	I��x���v^���	�-�W3&��n纇d����K��:
HA2)�8v��u�z���h?�ݽ&#���Y������"z�-�p�L��4��VDxN�p��(?�xr��g�J�z|���Dm��	}�!m�J�9Ӛ�1�Ϟ"����$V-����K@��>{��/
�=�<\B?�>��z��;x���ƄP�-^\Q�2�_��o�L�,\��#��V6�=��W�O�uk�������w�p�<��&~Ѭ�q�����.�B�wV
7f]�č�R!D� ���Y���v&��#�/�&��E�$Yt��"W��V}���>i����5v��S���~�/Q�XU%o<cL3[kK[�����^ 9]���3b��L-�-�kʄj��n'2���֑/��D&x�j<[��q�\vf=�a���^����J�`��ti�K��^�=>xJШ1B�	%��!��Sm	 XވY���܏�-���H��y�S�����`����p�{�l��i[�N��u���!�Dut�e�:f��w�0����y�w[�Ն�w�7�y
��� ��=�<;�p�ᑰ����b����O0�~�UV�fH-����z�u�b�;|��Q�Uk݈m]
�n�Zۊ㔑��"�yK<�\~�D��U:w�2I|��e�H���0x���z�,%x���p���9��J�C���K��%%���wa�=_N~��7�Q.�t꿍��fr���@�r��o�/(��!<3� K<g��M�L6"@F@��2����7 3G�wDc�������Hl!��b��7�� F�`˙��Cq�ǚ��y�q�o4bM̀XlxVHYEB    fa00    1500��I�I���=��J`�D�[�5��P3�Ԧ����6xy�������f���/[�MRp��a�u�r�</)�G�Q\����|�օ�p�'�����R���{E�����K=pb����-��Ym�&�v ߯�:OXT"�)�[vY�E	9�o@��4938�]�V�e}[*�4Zá��7G�H���S˙�5n�+	RvN��ט"����B��L}��j���N�;��K�7�,#l���?gv�'(o���&埿�W����O����8%6��D6�d��ٳ��ϊ�Ü�@N�9Q��0T�{N�z}�L�ym}f�Vͫ��7��X?�j��s������{�)z�".����W2��c���g��k��Q�� ǖ��8�j^D⤆�T���9�kZ�ٔ�;뎞g˼ �ϊ4i}��M�"ֳS<QQ#�l4�J=�/�a����
&F��"���g!������Z,��6o*���#g(��G)@90��P{Op2sZ
]ND.�ܷ����C�HFZ� i6ߐ�t�3x^��N�6�=	�I���$2�2����T�1� E�5�Cq���	�6��kX;l����H��;�i�$�[�+��&_�����yj?%�N{�o�6�M�%�e�)��q�o�k[�ʉ��m~�g����_�2S@��������Lw'��kTj����N�AGf��c��чvT�w'ob���]K���\.��vRI�ޢ;eqy��l�wwa��ztF�[���.�ե~܉��sm#q�����w�޵~c!��B�9��������~d�P�ne��B��)��("���0]L�*y�ۊ<�xZ��|_Ǻ5\=yrc~�j��N'���d:
:�n��(���$�?=����ߐw�����3Lj��	9T�%�p#$R���(�L� J#�)���XZ=�=�<N�G�Y�9埥d1�O�ֆSҳ��س��OL�	�i����Z�Ք44�*uH���om��=�O���5CtS=J��n�ڃ�),q�P�m҉ ���"A�%L����3��r ��D�ٗ�wq���t;��N��x-Ͽ·���-�G�ޞ�
�U�����-#�� �T������'�xO�����#FW�J"��vu���~F��Eې_R�|�h��I�V���>�Έ hJ}�@
�MԬ_���4��9���0L ��!���&}X��YR���{C�'�Q^R"�B�'�T'p񧍣b$��n�
�Ƨs'6c+
6��t�;�ʣ+3J��A�Kt�.��@B��ãX<���^�kȪ&��Af%�m�R��ts&�!��ܥ&�eh��hU�ͫࠧK���<����-��<���-���א�Eds�p�oZ'_M{V�5��V&�1���l��1�4f&�I�/U;�����܂ϧ���y2 
\&h��L�^��J�?���U�ʟk�0�:��P�${�rV���9[���_y�=(f��쿢?=8�V+ԟ��J����X�U29<QΧ��< VA�)�%�}.��
:�`�PW��R/����V@X*b�}|hfSr�r��2[�ԛf�(aI#�i�57g����Q�7@]2ŧc<Y��H�)�:���}��0��ʳ�i$�aC9J5�^d�|�@zG��T�g��с0�,�,�rX�&�'<��>��e�{�2��!��H�X]^�F�?ۮ����Ts�8lw`sa(-�����VF�E �9|��Տ�ݷ�r�s
�2>X ��_�꣫�v�Ҽ	�O���~#��lz��#98����)���J�n���I�r_X� �Ez[u�T��	�+؄t�����8��ӝ�W8���L���S���*r5�3�_�[G����B@��g�1'E�х-wB�LG�A�9K���j��c����mR��9V�'��?o
`K�oI�<)�,m�|��z$�����'�=��#[kq7�kl��cq�N6�I��u��j�~���E0b~|Ob-[�4�u�9I"�s�0A�M������آÕ��M:��sºtq�Aan��G�ސ�+	�������:�N�u��Z�z�-�NF���;ُX��+ǽ�����gm�!l��%a�ս���rK�[�'��'_��5�����s|ݏ�p�r>��� c*|�m�5Z!o��d^�g���� ,��$k�v6�LK�؊P ���vC�y�n8�G�5��;���.ŬFu^7gD��Wχ>r��S���w$�^�c/�u���9�Ļ�'zFa�j.�9��Rz�'P�F��I�ʕ���3(仞���#HJ�}�}?&����g� �5����@بz���K�jc�$�ѐ��Ϩxя-�Nn3~44��4��X�j�	�v���~'�'���nє�ڥCj�Ǯ]��4�:	adxcTы�ank�h;e(�G���L�V�\��v�ut(7��&��D��Un��r	��"�E�����\�(F��Ɗ�oO(;_2{64�9���|Z^	9���vc���z��&(5�5X��1�f�E8��l#�{7����v��.CX.iZJ�)8�Xk�*����� &&�0-��Y��]�ܛ�pzCo�¥5O.�l'ݣ�Ki�����E���d!�ІEE�n,5�E�ӵ�r���9��������z�Ʃ�\��E��L|�� j�G�i���3O����"v��1���ɧ���IH�A��C���T��!�X��M}=%6n�����I��f-�CR����|ܕ̉v�ꓽ&�[?��G"��y�4-��Ӗ�����i,8l �w�)�ς�:�G%�����}j�}��w�&\*m�=ٌ`i�ㄮ.UE��H�M�k�̂P�}~�K�<�i���ɞ�ۂ��R�mqf�]�Yi[����x ��!��i�@#Ol�ßS(��i���S4MKE�2j���\L�^u�~}&[��VX��v�n�{щ<�w���7�r6�rH���=�Tƾ��Vr��!�)�(�}��$I����"��[�P^��,�f�g��w�?��<��V q�Yӆ)��5��^�n�z�0h�([kR�M$����rF�x���
Q�
�Ƣ��Ao��l�Ҕd�4`��ܓ��d%�iE�]o�!�4y��)	8��3�SB.����;��Z�"%K�6SvX��$#r8��l1��4�c��fj|B�YƜ	�i@A�	��8 ����vf�R��J�wg��bK܈i!%c�l����:�R�� �i��H]<j�gGw�I��PXb��?�n�?}����{C9�����|h~��n�dM0&h�m��]+ҧ�p����
�u5���iX��O������4���,�c��=B����?��ty��Ut���P���x2��E�������t�[bVbV���#K�xt��@�I�3�w@#
��SV�B��G�(��aOks�HvC�}Y����-*�����t88P��I/�C��.��|Rk��&�,B�ۃs������Ac�:'�;���Շ'������:q ]����]�0
�\6Al�6В]�N"*L!%� K��j����Ȏ�4P��9�f����g`XsvLl,��t��'he1}d�JJ�s�d��쾘�:ƫ).���D��Hƥ.��P��%�z���0���k�ir�Wf�@���[�~8H���FtE��m��K��A���f�)���F_��[D��/%� �������<x�C!�j���z��	����x�Eh���3p���kmA@^e�:�:[��O����\����d+~?�L�Vc�Aw���#�́�yi���簲�s-ƣٳ'~wr*�kJ�^̴���G�e�-������u4<�g�Y�������*�ݏ�d��A7����pZ�s/n�p%��5C������q�i����Q��\���
�;�����T��͢ȡ�;SLM��Y��ݸJ�&'N����bWoS(�D�l^��i&S�L����Q�Ŷ��8`��yJ*�9W��>��_����8T��]�"�l�	�ѫ񾁄��ҧ+��V�S8l��ʿ� /���i��hu1J}��` ���˸xA����3K������{
���!�%�a�^X��H+�ٝ3,c���Q��LB���IY�*@�,o�]	z����J�ħy·yU�j�͒�:g�x���C�̩����~�u���,��ش<Rg��lnwm��3ʏ?��A��s�S�_��$SI�>(�ə����Z�0=�)$�RYF>�� @aKjf�0'������8��2�1ޑ	���D&��?�W�>�;�P�uf��� <Z�%Ӫ�"�!��)Ά������vu'�٬)�pG�0<�Oj}M�Ch��L�� y�=�i�V�6tր���}���E�)�t(X/�eH��h���\�_,4.��=vҞL3�&�,�ٳ��6�5tN�Tg1����+QA�?�{�|��m!
>�aa��<�]�A�5�~p�	��0�ŷ0p?��K~Ho>[�nc�2�LAj�eͳs�j�lr������k�BJ�?� �~�bE��ǯ�Y�8�K�wTXv��c��m��<n����q/�vc�h��B�`��~� B��C~Yɋ
�L�>��{���L'�t���2��i��j:�ɛ=l�_U���Tq滇�ux�����O��D��;0\�eT'�t��;�x�nU	��43��<����>1{�@�b�%I%�`�s�i��r�J4��ù_������T���D'���?�p�8�'%Q#6�OW�Sb���18�Gu��*WD����]v��YW���⋸~��9�n����J#zV��'��5z���%oRۧ�d��x��`���k��Ĭ Bx��2CpCOȗ��ɇ����ԫg�{P��%�P�mHA-a�h�P��ի��]T��[0�?��rH��Zh�a�w���ğJ{�/M�ὸP\H���5'��	{x���M&z�[�n���G�"do4�.���F%�����0qG��P#����yq!�V.�� U�*SPA��B_Ͱ�䞈��`�"��$3���G�H�c��j�8��7�࡚�s�W�	����_��భ��Jo��okVF�lx������'QR�޽�3>ߨ:��{^��F0&F�>Qf=[�����(KT��>����@|�����6pp�/Ϻ������D�z�I�$ z�Q]�w5�$�7v�4�߯*CH�9���ݱ����
e�у�\n�-� �4r	��ԅ΂�[���8��\��3�:<�b�,:P���9p�X�v9mz,��>�'�p�bO��=��W7>0v��G��,ˌ��IXlxVHYEB    fa00    16c0�%���� 	�uH����G���l{!����{h�ӻ���)D,����M_�E�_��MG{��R!�#h�s�0'��^����aq�'���P�:r�*6�ω��4���Pʻ�^֫6X!��u-�����E*��#��̀��q�q$M��_7�osM";�kg��H�&���S��@)�py�� ���](L�{M��uÓ֛����_�Ws z����?��ݻ�]Mvb:c`Ȳ��ާ)�E��6yTr^�:m���]o�7��-�6Se>�KIp���Z�Xh�H4Ur|/|����Գs��l���A��0ژ)�h:`�Y�@y��U��c:�%;11� �y^�D8pH��,_�X�\���Lc�jO�3iK�~�4�'[����!ö�8F�K�6��h���"��
U	���!�P�#����V}j!��5���Ŧ!����H��]��p�'D���*�,t��r�8�N�RN�*�9ƭ�Ο,#0HQ������]���P������o������Ш/�4��xsޏN�A%�,��1`T�����42{�4{f@��ly4���џ��,�LN�,�ݵ1�$P>�Wp):Ӵ0��,�7���A��b�kzq�3��.�D��'\�А������A�&|t��;����4��W��m������0�|Y�<��wkX������?(m�L�~����4��@'-Yc�4�
��"�E�i��ґz,M��ѝ�	����FaV[,��]l��&�
����.[�����Zh�P�b����o�D�n�#G���&F���T�h���ue�o�"�h����3ˈ]:t煰�����3#P��d_Q�y��?�ԛ���6���*��jX�30������� ��?iԸ�@���|��Ɉ�R�޲M���bJK�_�������<~��ЛV��7?9��	&�,��<�X���)hy����Z��N����)Ԭ���mAQ����@�-t����uh��T1��O�������������`H2s���T���9A�!q�@69C�W�'�{W�d<^i?$Tft���Of�����;�U�~��{1#\8.�m�c>��tф[�g\�)|q|K�t�'�L�d��?��\٭���ǔDOWC��5+���yɏ��%���J����B��Y�r�������]6z�U�%�zǪ��Ҋ��A[J��1j�8�~]&$D�b����4��8�(&�,�I�t?n ��>W��{���h�ث�Ϗ�9Z�p�S*�I��N��lR��_Xh��ŊO��+�Դ��ZW���\a��ݎfWI�eу�xS���9ܴف��4��:|��V�ї�BOw�s��0�g{�.�"L���8���$]U���OXN�i��T�W�����rd��nCƵ�xo�ys�_,Tgly)ٓ5k4?�GD�6|�V�a`�5�D5:P��#W�.Q�lu�����ۀ𑠤,��g�X+̢�OO�D��(y
�Arw������Ѫ�Ӊ)��XR�j���rw^E��>S%oϔ,u�!�3�+cd��t\���b6�=K�e;�Iฮ�8���t6�FT]�7 �6hp�9$���6<o�
�/���bW����O�fc/āN���Y�I������U�m��튢wɶ�����R��^��C��2���ʊ�:w#'�ۿ�^����	���'$?�r�S�<�^�{G`ls��B�
����\�O.�	ѩ*Go�(u��J��V��o�O��7�z����K�BϺ����*�p��,�S�U���F/�����'��;z������JP���[���
�&�y#	=P�j�������� B�UT��Q�NK���n�=�R*e���Ȇ�3��w[��{����m@��3Z��	Md��[P�Tt����w6c^s�
y���nL�\U��c�C��;C�/���9�=�H��=�T�b�0�|?j��p��h���U���3�p��w�h�Ku���M��y�0Dk�\�e���n(�d
�}�(��x+�=����p�r���w[�[i��0��S��ز��S��]q�<Sx��+g�>���Yf�����hk�."�y+�1����LŎ���T}<��f�f_�f���P�S�4�� �g��r>�	�+�b�D��yf����0(�p�t���U:E�;�0��a�wD8!p����)���x��/�t�"uR/D��^������)�i�M��ɺ��$4����ӋI�jT���}ê!ΜD8�P1)�����e��A���熄����)�J��{W����N���p噇�[��_�1{�W�l�����b1��WI�Z �e��خ�0gQ�dK4�؏�x����g�����5��Q�"���
��E}�*� c~f�(�w�`�D�,JӅ��k=���7n�_ ��� �G�h�1LFI�����5~�jC Ǎ}-[h��Yߝ�Z�|ՒP0�;pV�q�%47�,Lk��j�¬���1��`�v�zʉ�Y���;sdn��d���7 `d�NR2R�qB�t0���&E�"�U���1�`�QRo�x}x�&��	m�*B4������"[l�?>:A�W�A�Q;}�E��z�:M!�����$�e�ɶ��
���sx�C)w�_�c�o0F��C�UkJ����-�P+���ܦ@�9�2	]{@�]�Ya���XE�����w�8%��	��6L�H�_&7�o��!���D�T�����&�0 iݓk���!H[|鴛�eМv]�Q_��>��ªiA��/����nR�= '�aL�J��(4���Wٕ��b?A��G��7?�f�z�X�A�9�^�o�S�!��>g'����ӎ��W�2d0$�=>�[�L����?/Tۼ��Mn�@|6�,'�/n�Z9��Ƙ��k�Z��.�qm�2(���{L}��8��N����<r,��<�j��FOP������o��?���9r�����uIt�>?��4�ǧ��ؑƥ�p���j��`9�p���0��NY�~/H�}�0AM���I��Vʠswύf˼��U�m�ٹ�YH�����\��žJX CU�ʛ݇om�K�Bh��F���<4�O�Ì��]���U�*���9OG)[^�����$ɫ����./�氩����)ouB�������3�>@�q��W���h�nx� P�*0|�N��DX&=�9S��u=�X�U�*[��K���п8Z�>f�D���`6.o2f�{ڒ&��M<����J�o*^�I�����d�t'c��(�kk)�lT��*w'�ΌVB& ���>Ҷ�	,̔�p����O������)i���M�s��/�Xf�Gr���˩�:3������p��y X&}�Ӣ�?�K���x� l�|&*��x:Ӄ�~-�2��i]�Um#�nO�<I�V�o�o3pQ����e,@�`��۸}�i,�'�rQ:��5�sL�3fw���r4WS�9YW��=m��/H1����ԯ��d ���NK){�J�5��nM�z��V�t],��ťTp��x��s����,�
�Uz�Wg)���(���_�E��"���|'�ə�3�Vdg/Оo�{��Ui��d:�|[_1�G��&h��$I��Uؔ����st~��B.,]Ůt�kʌ�(�w�!S>bR�C�?H[�WM�Ĝ�+��M���b8Oی_9>�59�ߍ�|��1efh�{� 5�#����W�v[�_��Ec9���X�ˋ(#���;�"�5��y�R����N.��#]��}`λ���	����9�
Hπ��>5Mhk U�ǆ"���J9��Q�� K�
���M,�q,��(�D���gN�¨�I�/�sM[��a��F��Gg3���w�v8M��9~��O6��`�7�(���H^q��*�(�Nb�V�.k�5�e9^4`B@~�6�u�=��(����>1
t�l>�mր�Ӣ������g��v(�^���G{56c2�_g���\��v��K�s�D�� bJ��d �tF��,�~�c���6��`�Ų�)~�<�)3��/!����|������W��ΒZ�p��	�3؎�]�n�#49&KG��>3�M����F&��A����!�ͭufVq����z}^�4����L�Sy[O��%+�� a���/�m���w��Xʮ��c��H����	���| ̈́}3L�A~�z�}Ľ͉b�aaB�ų�4��>ë)�hH�þ��Y�9#;0�t�Ii�!^���u��d��&0�ޙZi���z ńtE{�&R�Osc�z��>�\yNN�n�+�H5"�c8܃k�E!��zes��ZQO�y�0b|�"��,%�~��&HCf%@CC�����o�����q�8\�K:�乆�^�=��D��T��핦-����,� �V��@.4��	�|$<`��j���|�?�҂�^z<��đe8�V���d_�@~6��ݜ5�jru� l=�Fj.�kwQ�	$ �>��;�-�d���w�	�������Tv��8Y�$�B��^["~/�s��(i{�`�,��{@��r����^�nV]�F�Ǉ���wcu�N����w����d;��5waĘR��[k��:��u�z$d��zI�GJ�қ��\u�5��o�%>�%"�&�$߰�2�h��D�qH�Ϥ�Q�?E�����l{]gL}���s��O�����4ߧ�Gu���lp�Ƹ����G<���~ �:��!O<>vrEܮ�l�;ɸ���<�x$g]I�"i����X	���^E�ڊ�h�����LX���<+�����睖�����?�+I�QW��I��7��O�� `�t�p�h_����x3#�kC��R�>�����t�����!�Ѭ!^��'�r�~M���������A.uJ2� �R[�������T�Q��4n���ͅ4&�OE-��4܇��`���a}4�+�C�O-��<�G�"����%#�_��t熤Z�Y�@��'��q>ͪdM˿//��6x�wO�B)��7��RQn�3���ĺ��sag�W��C�<�V��y+�y}4/)JZ{S��KEt@�tX�p�Xے��ݨ��
Z�(�'�e�;eZ�𮿡1��� �Lv�1j�s���<	xg��A�.��>:�,�H�Q�hdJ����@P-�@�^km	Q���w�Z�JZ]W�Q�6:Hb�I�x��9��Lc�����o�N���3�*T��!XU�p(��Y'��|�,�Mf?|,�:��BVH=� �P����SR��Ag�S�j�n�5$�a�;S�2/��]���% �e"Rh�wï�ە�"���IjT=u��r�k� ��:Zea,�`��C�+�`��'VV�C"�w%f���WhEdj;���Gj��~�ȉc*q&��q���c��_�;�G9<e%Z[�6�,".+\�ު4Tv����X��c��#�=������c���	a<e��<�3<=9��낵{V���/X�{3��iD�J 1���n��_S$��{7��`]��߲_q�-���	������)�Փ�`v��@��.ӍϳU ���#R�u���ν���B?&n��o�dW W��jȄ_�`���{42	]-�7c��t��3:r�Y���'�uk:w�[KEe\ٕ����Ӗp;zU���z��7w�pRlc9~�G�Q�C_5~���^2;Җ^�͈�>\�U;XlxVHYEB    fa00    1740ܷ$N8d!iL��I���i�b�nw�D�vl���ޣV�]է�&�č�v�ڠ�؁R5�H^b�����L��ff����^6�ct�Л�_V�̀mw2��y��"g�xC4;�b��k�};���I�Ԕ����$<��r��� 2�$�2A����q�����X �9TDO�R�6�"��e��}�]*�i��dN'T�h(�N�x\ȵ1Z������������0cpo� {V[�Ũ�(�n5/�]��~?e�����������6�4��q�ܕ9�9e����6"�?s�c���ęxF������ڳf�:�j{��5��b��#�I�T6�����D������7/9w�����6Rj�ul��~��F V���8�/��������DT�aT&�wO�ʻ�������l�{�^:� ��ƴ�
F�텸0���D�N-�������}�a���������}�W��w��W<Qm��;��*�P�c"��"�ػ����f���6��h�K=|�e'Qt����~��ɳz&\}�B��޹�/�b6&��z�2�8�/L��pD�|��G�K��m���~n)X��W�֘��
a�7�Ƀ��*E^��1 �k��K�(�p%�"��h�i����[U�]�ç��eě��V%Sj��!�����O�C�[�)��X�,-<��x�iQ6ow<��[��[#����q�嚖��\���d�8s>��S��f.�즥OC�M��g،55���=����o���J��{%�@F1eR-
-�2����<ݙ�P_�&���#!��0ċ�}���A��]�^)�$ئ�z�9g���U<��B��a���-�O`wL��nԣ#%�;uO�~1<}��m ł��TCla�_�����"���
�	\�z��1[�,͑i ?c���w�����9V�7�&XӲ$��W�O�ne�������v���##�����{��0z����N,g j�����~�}��,���0 �pK{Q�
�X��DWE�B�?_Ҭ�HD#5�i�/
]G9�Z{�Z�ȸ�*�*7ec��޾�f�_��ӵ@��*�ݍ�M���g���]Y����6T��U�aK�8� Y��~5�kȊ��{�jx��(B� ���(#Vpt�8�?a7��z%���sP�ի����x��2���Ġ�Pǡ��}���d0v��2��k�u�����uUS�w�Rr�^E��1�!i�u���tb����"�7��O�Y�:���ٿ_�S��>e�.�%����֪*�-���8��8�^����IcB����.~)�~���x.��Ot�/^�3V���߷́�_�g�i�r��d���~���f�����~��V�1�vo�=��,���s�G�D�P4̄̓*�M4a�@���qΰ�1rMw?c[w��u�Qm���f����(���'�a�/#���a���KW� *zv���o�˶��#���3�;�<Wq�>�<r���_����uN*E9.�l�gMÛK=nq/G?����T�	��
;n���p�	��_'0�FR��3ģj��������JhjP�x )Et�} �J��(��5��wf��D����Ce/s��L�dmg�a [�� �\G)4��w����gt�v�A��4:qe�oq���=�7$u�Cd�ʧ�P����x�P�WS�M[׎�����|E��}��Tf���qb���hE�<Y�>x����Ӝ���R��ϊІ�ҡ�&���6U�ј4h�Q[&��=L���w���'}���>g�V��V_�`J����Y����'�/�&П��[�ȠΉ�y�^���\ه��V�5lr�P/{���£u:]<�������
���p�j�X�$�D���<��"q��BW��L��j�G��C��f�hK���4��X�2�<��G¬�Q�L������2f(̯�`yjZYYl�m�5��qp�`u���O�MΨ�F�V�t�E��9݉�i����T]dQd��s9d߸T2����~�S�}�|lG����+1/��h,y�O.T��*�Agk�-�%�:�`�YSK �B���G)�!(wLe�>��&^��@�%�X��x]����[ⶆ1��6�9j� B�YJ!	z01�fc��`�2�yWת  ���AӚ7�m�wg�Cۜw[A��#���A�:�	�p`v����$\9��Ϝ$�s�}:���y�'��y��2�B��LbQ���$��6:_��y���k��U�~;*<�l�f��$�5��G�K���zuj������K����!uX�q诎F�y���yY����l����3	����Z��~�.�����w�[:`�M����W6��95k8��"z�XƋ�@��g�C@H+o6��J}U����ұ���%ʞM.O���5��ʐ=b�Q��5�%�"�h� ��o��>$y�8�Yq�Q �aP����|��nĄ��T������H!��u2��P)�GV;�t�K��i �_7��?�"ٜ1��Q~�lѺ
.O_9T���L��Mz�K>rYX)����pRv1O��s�6l��er�l�B���1\I[��Bܦԓ*�����]��!o�Gȟ~�߱�O~/��y��`�>��e�F@C���J��'����s�B@ąD�IG_��>wuk"ˬ�'[���4Z�+���7�oM�d��\�(|���$�}�������É��髁��ＥIȭ�V���������4�KC?���M2��W�r��DR��>�ie�c60,\ư`���b���&쫩�
�cV������Wo�a����1��{a�������Gt>�M���l�=�v���Ԗ�s�5���C��o��	��l I�f�_b�>t�K���w��0$������A6rcH;�.w��G�Ie9JRU��`M�k�={H���?G��z�����.��*s3�t��  g��h��,�R��V�b-2�Ħ��ǖ����U��Y���1?��-��mZ���G5&���ވ)c��E�.�(�/��S2��� \�hKP�������O�X�K�����O8�h��AQ�x-����OOi��{�=��C�W0�j����њ��9$x�08(R���[��ʟ�/��,4�3�D�F?�/~F����Jj�˳؏����y��W�ӯK�b�$ו�q��.q�����tIQĝ��-���Ph�nX��ݹ� }L�>���ڒ��r�Օ7W���v��]��JnH�>=�f'�uv��s��n+=� ��;,�)C�K��bY8{� K3�z� �6(%/��w5��*�����b�����@���=�<T밸R銨�C.g�;��J*�Y	������o�Y��1E0�Xh�/屘�ֱ��o������Y�8�d��~�����B��іb�1瑣�����z�*G��k��sRO��{�8 ���H��5̤���q�ğXi�(g�����i��\c�P����LV|�h%���,�[;�a��ƍUﶮ���|K�v� �3rDv�a��h�
�~t�~�)^��	{��e���=a��V.3�.4i�N=�w���I�{U]�A���	�ˀ���>��H�cm��|��HB ����{��t�&�@V�ϳ��Å�Ȳ[[�(�GHw��y����%�P���
B'o�����<@�b�:��N$��$_���"�Z�a�*���t�?HO��0t�� ��Q������o;*TI��[���rr~�L�&�d��hp ��W�u�D�7�mBRy�(�t����;Ly�&�!�vT��M���p���k���M�����g��ӛJv�y�����Ȕ��5���QA&�xIn9�dt��LO[��bǦ/Ӗ�z�g@o��lq;W� �Ux�o	����-ae�»����;�����s��Z>�[F��&ϊ�Lha����d�����0}nd�.J4
�fo��̠���ad�ޥ����q�X��u��Ի�&��lf��$����\�=x:Ƃ>3ӱY���H�G|뼑�$��g��}zH�_�s�T�Wފ�.����/�M4oiD�S6
�m�um��D\ˤ<-8���<[�����R�����J/��pYŽ/Fz��]z.ԆRԪ(�C��l�/FP�f�S�ye���mS���[d��*��7��'���7Apk�H��'K�tSq�ro�G}���e��@�U�[5��,��s���{N|-V<���Yv�mZ��궽=�$_d*�&(���!��ҰGKVc���R�U��а�5�(�*��y���%+ ??x>�:U�:'���ث�Z�PXC���UUw�����I�\%b�DS@�b��))ɳ.E�#I������YXmm�b~鉫���|6@����|=�J��}g$�p�����"8k�D?L�Y��>�Ǫ���-��p5�Mp��%����-�aaA���8u���6�nQ�o���g�/dx7���||��8h�,�dֶ�G���,�� [���lŅ13kS3ʆg�3�}�>r�T�,O��o�ŏ'�M�Ƞ����n�� i�3��,fh-���g;85H�!8]ъ�X���G�S)�`F 5g�p<��������J�� ؄�/�v�[�m�a��i�B�7���P��Y��wC�<���Y�=+�k���$�"<��x6T���rs%�%�"�}�*�,U`?H���R{]!��ބZ&��}n���m�I~8�
�x��w��*iv����آU.Ctg܂,<DC��&�1�$��)C���� n�_�@tT��3�u�,��]�/$���>4�&<V2�_ʰ�S/��;�%NU$7q&����%>��ٛ�Eń�������-d+V�Z,�B��17�IAI��(B�HB6fU���umཱ0\"/0d����q��ΜS��P�;��(cI�?݆�os�X�x(�F�V�eS���>��k/�KJ�?my��񡚣�!ď�����o��Iv]?NW�%�KJjy�2@��z�� �72��!�Y��������ŤR���$���G�f�Ϲ��;d����nl��橭+��ɧ���n7�f��.qת����V~�r>�����T�^�J`�:ֳe��Hk��:F�G�&GO��L�4��M}H� ��������ezqO���&�r����e�w}:�p�6n��{����Cy�sX�+]��1���;8]��3�l�w���_@�gBð���LrҬ+/){*�~���e_�QGry�Iw�HaG��>F��*1�+���m���N�����+Kl
]�:���.Tkw�����K.�8@��2|ig�.�Pg�bx�[�kJ+���vIa݀�'��+�nk��2�\����pp�2�_�>p���a���̰�0�f2��r���F�B)6_�R-JV�\ߦ��z�������S�uFi��$�\���9s��<��!��3/�ؘ���,�R���� �ź�ڬz�� ������N{}�$\#�l����r7��U����*���$@N�q!�fr8��ʷ{���w&�����Ԙ=��r��!���V��{p�G��n'r�_�����F�<~s�*�9�'R��b@�=���Ɗr��(����2ܦ��t�D����7G�XSO��� �����=f[� �<��0�k��7��8��_&�����%U|v�34�WL��g*h���L��ć�����Ҹ���|n���L����w�ﲀX&�c���U�8VG�Vd�� ���ԋ*�>�Cw6�SZ�J����9�F��O'�|��D�0��)�M00q�zH���)<c��:��͢��Z�{��XlxVHYEB    bf14     c60��� iޓ��O:�<��?��I��:�
��ct��̟5����
�?���m3��TY]�3��`�0�8M�i�ı�^�6�NZ�o�4��\��tm
C�gF$³�V�nuԶ0�9f+�W�C^�:{/?]�����H��h���nٺ#&��6��@�}uL�\�sU��uz�E n+ǨY���=��^��q�f�����"S#���=3v�Eo�s��q˨�l��z,������.kՍ��qR��\���n���23���Ex%����s�Fb��S�2�D�7�M
4#Ď��.�W�[SK ��K��o%-2O��U��=�3������?		�F1�n�aNJd���s=�F�چ�q�聨��6�К�:��˕A��ip�����#�/��7<s�}���j�LN�¢���p@��f�����Q��Q��6N��yR/�����,9)g��n3�$�#_>֌���{�d��c-;����t-c��i)�z�Yb+	T;𿱕D%���W�^�={.ًݝD\��e׀ڦ�w�<���!w��l�8�bK�$��Ԥ;T���q��l7��|m:N�{1�݉��B�x}#D�?��7( ���&?��};�LY�?x�ₕ�E���n�O�J�f	��3�����N1�Ȃ#�@Y�	�^C��W���qW�D2Kt�'��.������Pm5��u�)W]��ΐ�)�Ռ���9fhl#��t:}�w߯|��D��|)��5�t�4 M�!!�u���'�t8uW�Eħ�d8%KC#�h��Y��Ս�Q_2�����_q�\���pna�D
�`��ӳ�h�aZ9{�6J=U�a��[�$�s�P����K�IyH���f�\�t΋�#6A/��5O��&/�~�/�?_~Z�(]�d�@��7�Eg���q��Ú]��ȵ���+y0�? ���{9�H�T|v�Z@������OEx�+|�x_�t�X^�X]M��сӁ����g�P�h����kA+˨)����$Vˑ�����lA�-W*�H�B��C`pc��=�{��N�{� �-,�_`|�@����7�������17q��E��+o��2�3�_�k��2���q�;T���=���o{Q�[�z��0�'�zTt�3��pHd%�d�k� Bd�7CM}&�K�SD����^wr�g9�Д%�h�Ө^V�W��v�E'+�����]�6W�t�\Ժ��Ck��v��{�ԧ���r�A�l������2�D�����p����s |Qߣ��w���Gf���Tb?0�	h籂 I�I�l+�&��H�؄1Sq���kZ���4L�E��N$�I�N���к�׺c�\�%C�r��ڢ�����F��RA�����. uB��4�&߲��d6�F�X��܇CLok$��<3 �3
��E i��ԩc5�k* �j�����:��w��P�k8�Ų�7/�7�1s�X/�,��{3S�D�̺�)��(��5(x4i��p�F�B��s����e�2��샺�v���h�����˜���-��h·�~b�=�2(`����@���g�Eu�N�� *�����l��.N~5�C���u�V.�霂 (��	��Wf�o�>.�+=hQ�����.��}��@8�t�f�W�rݒf!lJ�D|��������ש��I����Ƹ�z<�����ckԩ�1�
@�����	��/��W_0�����I�e�u7=�������0�0���e}�ݛ�#qU������ʈ�P�V�o�)��X�&���k��><G4�	��\Jn[|l�F�)����*�G�!Ǵ�]�������b��Yk��ږ���v���V���c6A�&n���
-����j�vڪη�m�����Ec����n�J��Z�K^�����9bȵ��M��ݩ�܏<m�iڈ�$���	�m��B �"���niuez�%m�F=���y(6Jo���d�}�b	[3��7^�`;v�� ����^�}��!�/l��_ʛ�����D��<x������n2h]���3����@�?H|j��/}?b-o�Ĉ�3�����-��U��O'B�ߌm�<p7�ˢ:�\Ԏ�n��`���v���� XV"hj�WU�X��JG�RGbqi!Y���.��qg_)�7���b[�n���`s��u�ewcpN˹"@D�⎪��[<�A`'M�[�N��B��E���2�\:�w�0]A���Y����p�q~���f�������Nh%m���I=*�w�����m+l�ɛ�ѦX����8�ϴ�o��&JH��J��瞁N�\i����?�0��CpT�AW����I�������nM�̑r7Ҽ�F��	�sQ��ҜѢ����O��5� �	#Tn�_�Ŵ
1C�m���*��;`}����gŧ���Ce@�aq���M�9��R���55.�}_X�ק��:�ں.~�h0&��Qn����Y�v���+�@{�oy�2
�q�,�21an� j��p���3��:Z���@|������=`&D���bDƶ0�W����Pvޟ�u�3�W0���7)s6����x��C�W�XA���[�J$x��	�����_5�t��?>������y�
�D�
/z^�6���z|��Q�� *d�<�8 ޯ��t�����ю��U����f��g�;�tV�� ԣ�����4A&h���
�4���]�]�Z��8\����JLk�|����ȁ���)p-jc?�S倠eV���\��gp��1	
:O1=�
�V]�M � ��r��t�u�{O��P3ҼS�.��!C���Ã�''vv�*,+5{�~$��.h�)t�R�\��'�ɼ��=���g�J��b�o�H���"���CAX\<~�`<�Wx+Ğ���H2)�#�Y���<X�6�碕c�&�s�29S�~~c�V󀢓@񨂒܊���M����b8ŠM�4�QA�p8|x�+h��^�e�9�U��^E�aۍ~qRȜ�b�ݟ�,ϯ�M�n!E[�v�撯zq�$ᮆ/��������|M�[�XU�s�#O���)�1�n��W�c�xz��y"^�