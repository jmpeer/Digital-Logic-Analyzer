XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���vE�5��­�#<�HJˑ��Md�%K0���F{��d�{���PfB��=���{\pcå��4�����\b<˅�/�9R_'���_o��D�6Z�J��B�9�d[M�oo�� ro�����p�?��ߤ��6;�bRe|�G�l"
�I��!��V	I��:�{�U$R�B�Z�l�.Ȑ ��m�Gp`M\^�WQ� � t��Z����{����~��O��B!ܣ�s�������^���^�����a��"��������2*��Ǘe�@,��ns�rꇃU�"jW��~�u��FU��a"��J��3�n ��Y=�B	>4�0�!�/�˄ge�6�F.�p�[�'d/A�+-e�?n#²z���Ҏ�l#M��<FFe4�Z�W����� ��+�IД8"�4^�9Y����8=�/�H3���>;xm�w���U��u�v�#{� /���yP��"�쯞Q\ �M0kt�hY?Z`AS�_��{zwoo�]��� �\7'k�$;VD5�=�|Y2� � Ԃ0�����}M�J�,��X���z[8�p��ў��j��xt����\�&�b2�;栻���7)c8ܑ�L��7Gx�~����b]7��˥��%�{���UϜ~P��R��>-b�#8��&l>���� ��n]�<�9����O���l�����9�1�xG�������&�ר�cw�J��Z��R�B�\h���Hw�1M���DnX�}���;ɒ�*_%}�0!�>���Q��r���s7����_�4��Y^yXlxVHYEB    fa00    1950g�����7�S-b�>wg=DJٙ=P���m���26 ���-��Zc4!>�ɩ�b)7}��3C�����?h"�"��),���n�� F���R����P�Z���<��$�o�h�1�暳Dʺ���j,�=�)����m>s72ef"�����i��]̧������ 8�əoE�TxF�0_i�7^�8���o˾z֑��G6�8���6�Z��S�/!��YS�1��L����ƕ�*�OĬu#M/𙑎�W�
�Z(�p�,q� �U�.��d<ph����|;�:��N :�z���j+���p�ᖔb�,�6ڀp�t��� ����@�r[�26��5���m���(��M��r}e<Y��L%6�S�5���^�g� @�F�Xʅa<E@�����BK�iΒ���r� �*��#9�,�@㠭�
 �w�D:�)��T�_���������t]�3u��_�>wcbb�ɖ��n,=��x�ǂA����m�?k����櫄4��l�mC�Ĳ�?��q���yk1�S���9��]����`������gV�H�[b]�!�����O��0�XJ�d�mB���
GGO�0~L1�묬��y(��c[��B������DNx8���D�QB�C�A?�y�ih�^��c�yhd��mZ��Mt2�˚���Y�$���!E�]��Y0jyX��Ft��?L�}ϳH���Y�	��ۥtaFjG%떕�E��!,� :\�k8��
=l�L�a�>ݙJ�B��~]��j�_f*(���/�:���IU����N�P�E���y���Yr�"���PY����	�插�m�yL�����S��;���7���x_�{e���ܩ��-7�_偰� 교�kv���Mr*���֧���3�2���G։��=6�a�����V3f�{��gg1p����G����Me0�;����>��YDuu\���u���Oq�q{���*������
�[�R�b��hFW��0�p�>���i����ǁ���|)����I~´�yF5�`�K�{����y�U
	t�S5�KXR\�]8B^���Vʦ�?𬝯�H�o���'[B;��2%�W@�b��"�|o�6�Ze��ʲT�"���z��9jC��#L�������73K1@�����?xd	oE�Cn�]���~�4:�}:6��s7��j'��֭�LE�b��ф4��zj��2�n&�~��J���z�6C*)�R�SS���@�K�\�}�zف.�V7�M2��*��@�\��mEֱ�9W�+9Mi�ج@�����?c���������P_��Xk́i��Q�Ԛ��_UX�I��&L=N�Ė���;�;��v�\za�3)�2��Z�ԋDk���߼�Pjbh�aYX3��vF�@<pܻVD1���d�6H��r�B��o&9ۼ������*DNY@���N?1>;�~�>L�)�$��e��7�X0;��m���˽��>]�|��ߥ��҄K֑oͿ�͝�՗բA&v���)L��O����דl�UN6D	�����&���c�vjV�>؍�BIx���$Yr��+X�թk��*dv�����g"��yC"��Ω�m�&̨�A�e��踚W�\����,Y���6_�# ��}�5:Ų>9�r������5��Ɍ
Z�����+kXXw��D�A��֒��Sr�4��%e9[c"ʪ�ou���wx��UWmo̾���i�R�x8>�K'C��-����,�.�cѡ��(SC�����2E��"�z\��A���S��7��|̎#����ڏ�ν�������?�{1C'u\&ە�e,����I��*뱭Q]ScV��Y08��	�e��p'�p�_����#ȯ*�r)�R�0Q��Ƣ<�/+�H?���^) ���zؔ���.�vdA4����@�̧���SD4�p�5����fBL A�g�Q����`��6w�����(�Z�]3{���aYW�/���R๶����t_r�f9��dm�����w5���rhqފ�<TB61�߭��|�N����"#?��ʍm�s�����Y�A{<���?w�F�yߔ��,Wv�)r�,�ik�T�=j8B4��o���Q��YR,^�Q����Sh_�������A��_�L��� щ��	KݕD��>���M������\
�d;���Gr���6G#�ޔb����7ib}��)u��]QZP�z��c�M�y�wg��	W;��9�cZ�[��[�bǗ{.G�l�x��`�3�F�p����.O�V�n=`�@���>0�݇�7��%�L/��շ���+����8ɏ�"�a�b�"�X�vA��`�N���v���I���@��݉^c1�M|�PRzېU�������8g�@߻c/?#6�������5z���"���%hEj�d�?�QKפ+�Io׳�*	�2�l�m�ᚉe��h^�����:�,�)�G_p�,�v(Y��/!��"��v�kd��v���@�b˯�>���Ӂ��wg�쎉I�($q0������P1qW�i�F�l �����~�vOg��V4%��ɺ�(�R�!���d��J�A(��M�ǀ04��!��W�$���ݺ�Iz��������� ���R��	��o]���(j�{ڵ�3���\�!
C=���s�i��u�B|;��Q�ũ�l,��k~M�Ļ��x!���w�ʰW<
��� K��)l�JE��]� mXj~>Al6�ag� �@]�(B���O돡~zv��p	J���:\�߱'Ä�/����}V6��� $|�H��-ߎ����K��L?༄!��*�:�Ƨ�_wߩ%�.�yI�̭����j�"k���?	A����$5|�ө͢����Ǣ���!���=��G�W��yv����K�բ���T�b�Zh�z�y�J�և
ݒ(ޥX�8�ƨż��U����^j�g���i^6�X�����j��,�9 �� 6��Z�r��LX�%/l]�KىrWրw�u@]�p@��l�&�T��G*p�+
=�Pn,%x�E�nn x��5��]�)���9�
��D��1�RgOv`�؂5B���QU��͆�aZ�`J�"I�����jI_X~��8ϛQ�y*X�w�v\ʢծ���M+��"9�_���QF&X(g���f!m �8�+�YA**)N�����w�v}"$�W��W��}�8�X*�x�>'ү����a(�T*�JzxZ�:L����u܁s�H�����s5y�i��'���_ �o����Ug=˜i{�����%krJ�u�$���j�#x�N�Y�6��{Jߌm����Θ=J�:gj����c�� �lVx�tJ��.�ه㙮b�{#
�R�e[n�
59�hF�F�#�Qe{f2��L#2������x���O��tS�܈ic��s�ki����ӻU��)%�uU��R#�^����у��G��8Ė�19���Օ�%fpG=�zZ�<�)N��h3��N�A~<Ց"/�\s3�H'���(��_u�cO�r�^1�#x����P[��(#Y-\Գ��I�mW^������_��f��<� �V�v��6�r�U�E;���7ɓe_0�
is�g�e�B�3�5�ZPR5�C�X��
D��U�6*3�#׬�m�l�K�㑗���b��E�Ҙ5ل�j���@`��Q�5=�p��i*%�m@m
��{�����0ת��p��oԂ���_?!*�T�0�ե���-eW���������S��%J!kJ%��1�jD4��z�'� 6�W�V���Gr��5��OQ�fJAXa[�7b��ۯ/A#�!c����e0�E	g��DZ���KO �$�>���Q��T�r|��"؟�9�f�>UB��Df�Gp�NpY�o�:��q�H��u��f�\��T�V� �KR,�'O�:����'��Y{��rEI�~#�'0rԬ���M ��6�K��O�W��bى�Hг-Y��Ї�����V��W�x��ԗ����,�a��d��d(�C�x5I*^c��*���puǄ!s(��nr�l�L�b�>΢�A��vGN:��z[�؂�/���f�"��8�����-�}��]�C��4���a�HD:��b�q��)E!��5��^���6u^������ǈBԣ�OG����6*d'�ҿr\c��ƊO\���£Ǧ�=8���k.b��0Y�d�ji%���_�	����'�S��:�Y�Y���[k�|�"($�'�F��y���7Ї���5��a;�	}�ZI�E����a�}�ex*EI�.J[H!s������3�Q��*��~E�m[�k�~s�W_Z�s@������<�t2��Ki�U���ůE����\7�iY�~C���d֡T��R���r
i���W]=��T�����rT���|�b�`Or|2��0P���H�=�d�H���_����B��'lT�Q�O!�_�
�c<#bQ�;)���	��@�J2���
_ui�k��т�@6��M�'���&*��� �&Fsy�2~V:�RJ�U��2��b �ϿFlx��n�B�A�/FC�����d�>+]ed�>ծN�_���[�z��B�|W����@G,,���mj]>��!�<�%��N��x"o� h4��@�@C2�*<w�V�:�v�*RЈ���Ŗ�(�z	�5�{4Tġ32�L�,��hV)j��2$7�����_������V�쐔�����uP�[�T<����e�AKYm�Ic&3e{�����"�S^EQ�c���+El������(��D%��e�c��v��˺�(4�E��/tEV@��<��qo����)08GĆ	��������_�l���P��U5�|fn�`Y6��HԜuW� ��^�Qѱ�����߱a�%1���P�\ɸs.�!�/U;�`�|ٓ�J?�*���/�ϊa���!�'Qh=E�'�"wϒ( �5e��H��8�m|�~\�D�3%����j�j6�5s���b6��:�$=���ed9���R��y� �yR��m�@��F ��'S/\	�����+\t���0C���aȳ|S�!�J�i�H<�����-�G��5/)���p��2JTPD��nY��=BqP=ɣ&�e�W�3��L�s�P��|Ǭ0i�����BR6yHҶg��}Wf6onZo��24yl��Y����F �~�-Q5���Y��R�?����q��u���yOUx?�ǃ�0���RYά�f��� k@��DC��YJ����5O�Rm�H��0.݂hGm�M(@�\�K5�Wn��u@#���Ab�����$��ņ�\���Ҕ��+���Ɗm��p�R��m_�x?�j�zB�j��6b�`��xîp�`�&���-ά���(o�?�����OʢuX�M��Y�(z4�H���c��6�=��3E q���@+	��Q�o�
���~s~�����YA��lEA���md���r?��b���c����)Ԩk�>�>	���a�2�4</}wW܀k�		�����ެ�J��;3ncd��`����6�e��(}�-���@�����36YfP�˵X�W�M;�|듄�B����DA�����}+���7Y,Z�CRb�@2�X�%}`-^HAם���.6��֟�u������o�G�d�h��"(��joӽL2TTj'�K�s IX#��R^łߘ�99c�~*�Q��k#fJ�h\.γ6v�}�*�`G�=��jv� >�_Y"�&�~7]�҄
o�Q'b������a�aB�$z*{��E�b�`As7i*ݞ����H���j�a�K[d���$^��A���ךJ�g�9r( l�KS����}��t�y}�+Wx�0t9M��FL�^�0;R�Cq ��:�#	�'�6����'����^P�����#�R�[jd��[��`���q2c��B�r�a|�"ct�^o�7=�
/XtF�<�1���A�\��`��}Q��de�D�d&,I"�Q0�Y��$�ALM'+��C<��K �u�N�D3Q�V�6��N�2�>xí�-�N\��l��8-��_�Ƹ� ��#�9E%C�`
�ϕ}�$����/2�[��	�P��\!�U9�����ߡ6����.:�t/-K(�sY끖�@;��śր�}�+e�^��U�5�t�����^O�K������T������t"������a�����������VN,p������i���� ����f��3XlxVHYEB    fa00     700vR$��(m����l���G�P��{KFT����?@9���"5�\����1���Ųy:��ܨP6@}��lUmŏQ�����ﴰ&ϓ�S�f�s�e�.yt?z.���WӲ��A�^w4������t.��^J��(�����L5�`��>���	��5�o�'в�7U�=�P��첳��I�qX-58�<��0�l���U�jkOܣR��7N?�8�SZ�,�6��b�W/�(����W/s���k�`d��F��HL��lm:��?����d�~����D�������z��$�	�k#灃t�^�H���M�B(�;2���(��)P��R�k��V�LP��i�8�$���EK�$Ѿ�Ä�R���Lj��S�҆y0"�iQ�`5J��\,��4��b��"�+H�,���3�xM���$� �X0���A�f|L����b���(}9�Z��S������*�ϡiC���.0��xiD��,%��xew/J��O�o�H`�RB|B�a���J��3Y�]D[� ��v~Z�����^p;�F�/=�O��G^���B$�14J�/�O�]Y��"l��n-�Ⱦ��d� ��1����¢�����q��Y�M �1��QɫpdX�>���^��3)�!�G�yl�?F�vi�+4��K1�Z��	7�D\�������Q���G����ߕo-j6�	%
�7�_jm��	�n:Io�A�E+'����
���y����{L�6�Ñ�>V�j�3��?Wuj�0��G�Qy��>�U�T���e���_*�G	1k�TDj|�Y�	D~>A�b~(���a��^��{��X���aw��Sq�B9�^5�_�G�j�y�������	1i�Ǒaf/�����F�mu.T��E?ZU����%�]��=LW��X(�á5�╙"���A����IP��sV��] ˝����)��'���M�t�.=x��a����.I�k���"�3��1�E �粣~��tRbŴ�m?c/8U����8Տ�	i��3�߽�#<me*F$��J�<�C��"�vaE����Z�g+�Qʍ� >���؋䂆�J�X,C�r̹Ii�%)�rª���Ɨ�կO�E�.[0V�G^�'�_ �V�5�C�ʄ����1� �C����_��$Da+W���-C��˼X�Q-=.0?"
�;�8�Ӷ@��(�u���Muq�~j�+7Yj��/����x�?3II�J�M��C�:����_�]G77��K���/��6��m}���Q"+�p���)YV��%}cVK��E�v/u�:��e���	��0
@���m�0D��' ���&^jŞ���d{�	�S�)�zʝ�(+	��QWn�؍��R'b*�r���B�M(�C��ƅ~fOAӇ7+6�}|�^F����]����ʳ�S����o+�ؚ#�$��?��P�}�}�E��Dhl�P�E�9�D�S�/ݜό=ǒ{y]�r;�B��m�@1�����7�)stGA��3���t���j�C�#�qŗ���Fb�e=Q@0�o[	Hzacܿ 9�2�0��®}1�t\�[�<�
�G�������U���~f�[�q�[���>���aI���+��x|����p���rپ�2�Pb��۶^Vc�$�����ɥtE���M����41����aYf�'��Ĵ�
m]߬�����m10�^�1�����Sv�(o�ԃ`��� �ri�^��r�	պ�1т&
�%��/a��!R�����x45U�Y�F`����J�K_=���	��WB���ZG �c��XlxVHYEB    77da     a60"ٙ���ʙ���� ���2�I[dXk���R��IJ�9a�O�V�FT����ca6�=��З��P#�N�	i���zm�k�PL�PcF�A��:2��de��K��\fa�}(�fH�F�d���K	pdΈ�)��gl���U���l�$953�����$�~7�=@�x;Y��{�]���u��t܉j;*��x��Dd ۧ\��fb1:�<c: ��ɀ�7�/R>�)�XI�_��1h�J�UMƷ����|D2��ǜ_{��әy�c��`<��9�����(˄����W[g�$f)��H�d���D����� ���)� tJ���	A��+��/5f��H�`�����۩f4o�ug���8P��x�if�F+�bT�wΥ�2����i���g��P����e���6$���D�D���g��UYl=1[!��d���@����vs�󕧭���I�u��k����w͕Qar��J�� ��e$�0f�b�.N�7�Ҽ��������ͪ���qn��!�$8���]�p����	�	��(��-^G�09U5�03����_}y=T��{9 �"yt. �+��=Y|�^�~,%��Y��r�p��%��a�2w	��z�
m2}�B����b�y)ꑵ6�R�:����:Ỉ�����ʦnҖ|����r�;��M�Y9Wl�b�c y��9���R�|�`�</,$K���y�4g'�����.�Q����_���� @�n�+�����V��>�Ifdq^T<�G>����ɉY+$��$�O{���x����8'p��p�|��;�ݸ���w�n$�7Pb�#X��1U���_�(�L�
��N���N�9��Cm�d���} �g���<wq�e<t��=�g�L��AmEy�}������&y�ńC���]��b �Y�o��zq��`��XdWi	�������h�S��Æ��h���/��o�آ��-ޚÒ�'�9��J�g=�c�eEbĖ����GK�E<����V��s����G؁��EhE������D1,S+0w=�*H�9�������N�P�"Z�����9�@�Cڸ7�	�^���ou
v�
�ЈXd�7䬹���^G�M��'tu�^�z�BX����쓂��d^��M]�P�&��N5C�VP4���.�B�v�1�;7j� ��kLQ�m��Gi(g� ���V˷}������'�� �_/���ϰsD���G�k����lur���N��_~�*�h��o��q����5[��=i�=����ZR(R�w;�ম[�
���ю"B��/  H�d�sb��s8�sJ�l����4��&݀ya��$+�F�:")˽���`�� Ţ�}�K��wK$n�{��(0���*-����Ō��̱E�4t��o�Z�b�\n�� vPcnh�	�	��Ƥd 
�=t�3r����ɲSPM�is�i����!�{\�-UO�<Ii>��?� �Ta��}3QTik�L��V���|xXft���pU$��X0r����ì�ʤ.�@\] ���S%=���+�8������޿�T�x���S���fU�+>�d	UN��)�ҹ�`����V�7X�w�K�H������atv~L`:Ҥ��2�7E�F3�	�����C�	@�)(��L���:��3�c�_��D�v~�=���>S=�{�1��m�X��7U��e*uGKۮ+��J)/R��5�]��,�`Su1��� �'�gJ�ż[7�������%��mH�z	�-@�A@G!:WQD�@'��j��Q��(�_�qwr+��l�S��XBq�] `�|,
���Cr:GAYgD�I^m���U�Y�{��	x5>����2d�:W�aߥ�cD�%1�2Ez��%^Y�η-a��Oq�6_��K���2p#���b�R5~��q:���������v��OC�94�T�Ob|�Ǡ7�B:�o]H
�>��m����?��Hv�*��<��X*�����TX\����(Wm�T4Mz��[mL+~����Z2���KG���dڰt<p;!�I�S�V-a�Ns"����
~���\�B,u�
}b��(���8��+E|�"�Ť����E�;x�Z8<��i9��x����ⳛn\*?�̎�-�~���H{)sJ���*?���*�6�
F�F�I����S	`�ia1
{y�����u��M�Yâ1\��yi��U\Z�s�M���h��ӄڼw�),U�A�k�1�P�p�}G �����F����ONvɟ��x�:�G:n-�t��E8�ʤ8sQ="�;�ʅE"Փxv���W�U���{��S�8��zs~p�5'���^]��4��v���K�x�e�k;K��Q�sOi��,5�����Ã簂:5^��FV�p���SG.����ܨ!��V���7�t�����u��ƃ|$B��hDw;�Bx��	*�_�K�ȵ�oӞY����d�/R�!q*��=U�$�وul�ng�=	�B��4vS4�MW���H� �/qG9��B0b�ޏW� �����ga���/��3�sǼ�Wə�d�"�Ҕ�