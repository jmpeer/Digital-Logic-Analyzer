XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����~�U����N��Y�T�Y�j��Ȍ��=Բ����*���N�	{ܙ�]}U�k�5��W��Z)Ь�ZE����T^���+��sz�-�3#��+�XS2��4n�Al%�y��엓:�qv�%�;N��<6��Ѻ����,��fql	q�V!r���x${�-2��k#�&��Ϯ5y(#mF�t�2Ì-�U��N�����<i[:�n�c���m������;�w�Cϧ�)ȦVi�z�Z|��-c5���P���P��_��s���߶F*b����?r{1�>xy S%�gnz�l��L���'y�ET�mMW�������D���F��pA24{l`SJ|aI�Ik�}��/WH�E	��P���5?cy�����;���>'�H3���Um܂������8��G{��qc����X�Ե�q�(�N��h�ߟ�gA�0�E����F��O �f�^����%|.�3]v�Í~�x�]G&.����$h 3L�4����[�g�����અ��-h�]��_�õUl853���7�K�� �� Z�l�%�o>Xv�_	�Kd[W�AYV%#�)�_YH�z�n?����g���O���*fЕn�y�~�?#��D@�B�sa����)JX�}"V�㏌J�u���p_�|����Q��-ǚ��_UR���
f�X�K�Sd��R=��7	S/rKLʿ�ӝ}]I���½_CÄv-�a\8�d��Tؗ�9|�m3�����I��|&@���6�A>8��!XlxVHYEB    2e55     b00����3��(|e��$
���0�	E�)�jN\��5Ѱ�jRg���d"�pE�2�S��Z��n�"
�z.�*ok�J��/��O�cu>\3�ֶ����ǯ��d:V?�r��9@h��?���<�ڮ�qԵ5M�7�l��f��s�;l�2�eA�e�*��Vn��H
q|��f��Ϭ���`5X��6�W�������U�o�ue\�G��v>:BP�Z>Ҋ��� ��Q%��I}�������Q��=U����Y�#��3i�c���[�ћ���@M�~�Β��Ѯ7��vQ�LKr;ͯ�ڦ�ME���ò?��.y�A�WF�3��A�t��XX[\��,=K_->�)� �+�7)g!l]���W�ub���
sD�`��뾭?��fT3_�Wq��yă�/���Ũe�-|0�U���-:(��<�n�h�Z�PAi�Opd�,.��i�S��'hN�d�5�������y�}�0�c�{���Yxu�$`i����h�	��~+�흏8ܞ�s�X��wo�)�
�e�_A6�Z���{���Sx��Ak����AK���"��"0�=WcT��y����%ZH�G��)K����W�e�i,H g���h�u������K�!HKV�W�1���8Cy�z�����N�Q��tl�0ķr`��6�Uo�@�0v}�`��X��\k�����9���TJ˵�a�+#��ϱF�]����;ܔi'G(+���bT�U���:U�@ͺ�C���(��{u������t����mg�8O�Y���{jP�w�9P��^���H^3��̱���r#}����m�x�ȯ�bo@������x��}������1�,^�}6o��79�	P	�&ٻ#OxO'%��,f�r�X	��j�U5�1L�E±_�޺�,g2�._cm)V��y��B��|�_:���~��%m��������V�i��Цh����:b��G5R^��f ll��bh~@��oX��JfK��mV������LR_8!����F���mÊ����ue�}=j=>����mLy�i�E�U��������]S��]]�Ti�r=s��χP�zV���r�ׂ}��^�l��4[����[ (�+���i��.,�?g�������> 9��"
��ړ��<�7,A�7����"���<�m��vFef��bV����K�B��Ԇ�Vs���JY�
*�}�Zlӱ��R�ݬ�5���$\�&��G��O�&�x$V�>��aC��>Kع�*sN,�>�Ę��%�y���c����#�Z���Jk4*����U7���޴s3�ⵙ]%���~�z.D���D�+kW��,k{=�=�r�T��@
I����6�[����0XQ>~�ߪF����uwh�%���z�-*,�D�l����ր����ΚsD%��L5�[����h���k��h~�i��u|�C�{'�c�t���/d�EQ�g�}<-0[?R֗�.7�8��D�J
0�v=�<��J����Lg��̈́n�<�l�����6+��X�vJ񒯉�b���˰�xS1��Q�Q�/��h��R�q�������/$ٗ���N�[;������U4�����n�So��#�&)�A'�'��1$V'�u�o��*��Iݪ~�^Cs�8ϱ >ĺ_k�z��m�.3����/��V��d+M�ȻM��˸��е�z/���?�����M�\����HϢ۳}C�(:z'3���p�R䛖2S�6��K���s�Rʥ�GL��� 2 ,��i�+���YƗ���P/�|�.I��A�@=�O�� ���ɉ����B�Jʂ��`-��og**a��X��6���0�
:/��G�;(��.��b�Z���˂#U�=��i�|�����������az�L�^���|fE^`�^ߗ�� �A�L��[����̪z2�;Jn`Y�%e�S��N�Z�z��#T�fI��z�T�OI)	����; �$��'��U��B�1��T��p���奈*6���]�*σ"��Zl�)���~/��Tu�s�C&)���C/'V5�( �y.���倆#��Tt=<�yS�r_)[��{q��c-��>P���`Sp��� K��a��������`z�6k���fG�e/��5�ۗ��Tq�"�v谅�;��q�X�j��%B�<ʝ��|Q7?��>�eP`ËZC��s[~;9q��އ�G�=�8�mWص�WZ2��P�5~�wbɹ�a�k����9��g~�']�N�|�'?��]�
x	�6�H� �.@60쑢02�x[����L
�#�,��J�J�uG玲DR��0S�#+e���N�ү�[+!7�7��E�h�/�	v,��sr=c=��B6���`˛6������G��?��j*�e..c^��R-4�t�S�=Ixڝm%_�.O�ON�����F��H�E���V)H<  ��������a'О
��^�^��1����ɋ{��^�H: �]����������1�&ѫ�&'�����,��e�\����k��$A�K9Z��v�M���Z6�_��������Km�X��p�oX�J���������\2�/,
��M%��!���5�%ty�ɕ:b��+L�<w��Z��/�$XRzV:�eZ#@8�aMiM=ƿ��,Ş�kb0�(��!.��ĥ|�Ĩ���'�����Q�G��%�����ܣ7
��ɺt�U4�of$�mHo���1�螒eh �+�e!�
E��=7����|����bB5����