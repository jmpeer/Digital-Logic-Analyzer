XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����Y�I�(��*N�K;��!�8N"&wȶ� т�zl9:�|��X�9�ai픒F��愴,��N}:^E%�����u�N����X�=ϗ�$Z	U�T��6�{���{1���ɨ��է��Y�ZlC[�������C���f�V%�+��T�ALf�;�٫m?ש��1Ì!9����ԕW ���D�R=�_[��t�NݧCIЄF����I�zR�5�i@�ǲ l�IY��2ۙ�aXR�6��h�����������������T�9�K�@C�2�M�Ȼ�b�W�
�gu�b�'��Y��H߿9E�z�;��
�K�����O�㜇
���Nu�z��ݭ����M����7ؗ ;�;4t�6Ĝ �B��^�=�F�Y�&H�˨�a��^\�D����W�(*�l� sk�b��}x���2\���_z�Y��O:31�����-�?e����[�v��ki4c����H	�p�J)�V"�nQD�T����ѱ�[�`��
 �}�����(@lL�1R����^��$<¿�z�ƕ�O;Jx���d�4��߆bL��7. x%�P�t6�.�h�{)���������a:�GE�ZW˓ARNܞ�\�T���}W��Q?I��w7�$ Sa�RPA,z���hR����B�1H���%�a1b��nHf���Gb�����X_�?{��1!V�6=�AtU���|d�_���`��bi���8d3'v�Ֆ&�!Ⱥ���<ص%���6#XlxVHYEB    fa00    2910Ht)�D�
;���Y>Y&�ØcǇ�m� H��4ˌ�*F=�M�m����h&\\�>��I�B�MOB�	eU?fb�mJ���Z�n�բ�;����i�q����m�r����)�%ȥ����#sB�+{�q�>ʉ ���v*r*�W颫|�i}�����YcC9������xX��u�4��U��Dv3euK`'������j�16d�gN�.dG_�<(�o�i��6�g�� 6����յ����{��V
���.�B)]y�������r�q��0�5zR��.wby��,�+ah�{�x�?l��cY���#�����0���\fv��UW*��U������>~eh�M�=�_�*`]��k+V��ax�Th����G�E��S6��@5Y�9�P(-���߼ ]�V���]���_�ϸY� �$�,nS���yMn2�����_�������C��O����Xd ۵0۝�`mG8�	�0��(xW߂'^�y�寡ر�������J(��I���)��7ES�V"�{usq?_x�`R,�d��HA~�2o:��'VaG�y܄\U�*��Be����D��V3N���-���
��hr�^���}O#<��xd�}?���F�3'V�{��ӫ��S.�XS����\f�O��/�N,� GaY��2s}x 0T�sO����X%�R6Gj\�Y��hP��EB裙��tO�3�YBh|�Ɏ��J-����hVx��Rʬ�@�R��q�($Z����l��T�y�� ��et��.��Ŝ	��I�R�<j�X�Q��o�@gya�N.uiđ-��d!r*�C�r&��H�/-E�w  H`^�Ag��wr��lK�U�q��J���S���s��V���_O�U�|y`B���[�(����OV����H�
G�344�=�Ǿ4F�<�1��R	�R���}�?F�
v�nZ
k�T�qA �ز��%�ٔ�@��R��S�u)��h�p��P{��a,���V�{>v6E�Mp�	G����Y%9�M]�اB�alrM�M8�_4�nF�k�tV*���=������j@6�%
�fkY|�|�H8��[�����Gw��XOm"�����B�.�(<?$,����:
	��Aʅߐ".���$i�ɓ�6KJ�ҹZ訠;��黅33X��D(��B$������Y���fjh����ʲ}�$������4���|��^{~���!`�0H4� iD�!��m� q_E:�~lX�>@4M��|�����(��X(<�AM]����bz�����u�q�Ӹ�e6v	W�ĭ�d,��B��C_t�Y��"���L���,f
�70��C��)�(3�r��]KZ{h�>�RΚ�����˿�Vu0�]�q���$��RU���7�)f>_������$����sO��Mr�)ۂ�`+��,�޹j���Ey..2Eں�֨\��Qvh�/sf9�{���+��)V���Z[&z�Tnm�q��Y���U��x��Ծ.ٜ��Âs&яPS���(�Z̈�/�Ė͂�E�D�Ӧ��=��a�^a���D(�#m�ž�Mw���k��a�-���9=V��;�8�y>rn(����3�նC�*l?�4Ml�3)�;��gU�8�8.��N���̹O`�Z7A�$i@�1�`_xׂ�U��=�S+�-��)�����<�
p	�2���oc��#�b�A{�6f�xh��i����ό׳-��q甅��ɕ��)QA�#q����8�M��b�ɿ�Ҫ ��͞K�d����-kW)ux��t��28.�m��5~u�܂��0'$���K�	9%�}a[ɢN�w����M�z ���;��b����}�Z�!Z.!�a�.�d;�����P�,@�p0���Q�������z�����ۈ~���4t�H�a�_¨�Y>�oTX��)�M�S������B��E`L>�U �rHSS*���\�~\����+$y�Z�x}��^!]q��p��ٝլD_�Wtcy����oF�0���<i�Dg��M�{��C����N�A��d�O:LT�>�d;xv��y+��+����m��<��U����PZ�i��-Q�E��uA/=����_��Ȫ�8�T��G��v�n���˩����j�_���f�yvG	�R��@��������Nρ߹�K'������JIc���
��e(�:��%�*2�Z8�3�7_1:��ɂ��T��`�L��k�n<�@7�zL����!��|����/�c���O.�:���bƠ�[���|w��>��?]��OuoצZ�L��}�36b�R5k�h���f��hJ�Li��4�9���&(��-��ۍ�4���ﲠ~	�p���欨�Ǽ�|� �,7�D¼N�������\���� 2��O\-����r%�<2�� �_�S߈z{}��n��������?��sy��ѩ��L qą�a��U���#�Q+j꣤�d�#8{WT���=2L%��P�vᙒv�C}_󍊨W#�ؒ���k~�a�i!9�V�[A��˱�B��m:�J�80�b6���F��\�;8����A�*1���W���Ņz=_:��O�#M��!&W�W��e̬y,IRZh����8�h�8I��Ul'yv^��ո���i?�v�\|s�n��
J�Ͻ�n!M?:
��a]@ OU�5Bo=]��W.0��glƾ=X����&X��NdA!3�F|$Wo����^��.�#��'i1D|�$����c�kf�(gJe)^�[A�n슬p8������s�������>��E�ǓNr/22gJ��X�S���Q`��HJiSJ��=�qb�ڄr�jJ�����̏�`/�Z.c*T�����=_��G�-i}�f���/�!�w�����Qb�V�~Gpߊp�8�����^�a�="�VX�M��rf�C�ؚa��W�~k��F��3י��+�R*}|v��3��'Zc���Ò��z��+O��%�~3�@.��I͸�$�?�BQ2�s $���Y�_�JYX\MK��H*���"�(3�j����+�8 V�Wh?���I���N;�����Kw�h��I��}�u�,*|����Jx���/A=d��_6�����io�A<�}R�G¨����]_���g�61V���K Uld"�w��W�lZ�2�Pt?�m�߄�X�M�u.7˕�4�-���J�
f�ȥ�05���`����,ʍ�L�߽�ӷ��vK����g��y�*sbm��r�ԭ[<~�FW-�*Jm�M��&�)>(��3��X����^A�c~�^�ffs�c��|4�xǷRy���N��H�H)���R�x$���A���%�(����@m��Z���:G�Q\6��z@Z+H����i�c06�@�c(V�&���ܷB��5�����or�)nHZ�uMs����]HhH���I�R�m�)�(h���٧q9��bC�����0pq2\l�[X�� eH}�S|��	+�*V�r���⍳@z,��F������:��5��25YD_�A���m3�������Z6L.Na�h	�i��-�Sj��IR�éw�{@xn�+
��#�1�����<�jI�֔�c���x%��H*]�B(k6�;�𺌌��{�����_@�܆��7]a(.E�b�Һ�Ï6F��g�X�hݔcm",�t!Zz�����g�V�.�R�9��ִ*���ڱH5�33C�����z zi3*��K��^�{#@��[))�'�^��q��������gK���~W���z�M�X�w�o����Dř٨ւ��a�x��h� X껯��ڤ�ЧǶ�39��(�[�T����oٽeY0��I[j��Q����s����%#�*�}��Yֹ�j��=�<�=]�P�v��Q�	��ZQh��gV��-���t5������k��h���7OB�~��������E QgS�����h�:�^V2ݤ0ꨥ�縘�1��S>�n�,��6q�$��Ҩ�M�6�d��(����ѫ��#2��樇�=b�?w4ЕΛQH�>�{A��])�G��R�?f��Z�@O��aTY%��%�>O��yՆ��MH+�<=�ۖ`���6�C�=���-��ȉ��n�/��eM(��U��#�u�B~�;�.X�#hp��?�������l���Ҝ����n�.o����Ƥ�U����<����ӒL�rMt˧��;W*���D��+�����F�P,cQ�������iІ�:��8m�+��o��y����t~��A&J�K*y�g;2�Q�0�
G�����V-S�{e�������0���������f7��GZ�A�>����10 mq0�;�l����z���<���)���܎���O�֨�ǐ�7t��äUwci��EB�b.�*��3=����P��׬�0�~�#V~�P���ʑ���2�dʻ#`��nF�����O���Yc��5z��D����6g�p�����^������0)����9M*����3å���Ҳ���2����=�?�nK	�-�*�\�A����E�-L��n�Zb�Ɔ,��
`�|��D0M�e[ø��� =0 �D�5�ޚ �å ~�P�e��bR_�v�Bخ�B�a�7�:m�{ �~;<�5n`MD�0ק�������Lv:�u��W\t�y^!�����s}Mj�HYEh�($�:'� �c�1R@�8���b`l�X����������T�(Q��p ����5�G
�X*�W��'Dd�E?�\[90Ǆ*O(#���0�(��BR����u/���k8����jҵ��_x��I�T3*/�vi�|
��i�x�����ec��R�iA�0���=�dS6M�sM�R �h80oq�x���7,�]���>���\��G�1����jhw��L�ϣ�U��'ʒ,A�$n V�*|*7@���J�dq�Ì�lJ ��C�A��`��aS�m�n���@�)�pYof��^Cm���+1`�v�V��z���/�;$g��ⶆx+�&b�z��f,f�ni��w���V9A������d=�s�T��V�Ra8�v"8�X
+��b�Y&���bO�>>d����Z� �p�  �s��[7C��ݽ 3k<�+5�t���7�� tѡ=1��ޡb���%����E�I�܇��f�k-V$k�$�k͈3#Z�e����d0Ffww3�CWf#����M���8	z�A�\
RR��I��щ5kR��Z�ۚ���1����Mf�8C�t�ˋ-}F`d�*Ġ��5+P����C|�9���0��=�� ����Pj!5F+��H��ZP;���ń��^���l��)f��9q�l��l��j� ��=�m�H8+�`~$��i@챠t.�-��]���4SX=�m+\�P�U���f��ԝ)>V�x�L��Ѧ,!�_"%�l�w8�n��>�����>bq��i)q���X�4U�C��P�I�E��O,"�H�b}�e]�t��1��mZrC���bL�i�?	�|Z�Pa��IrM;��R�j�;�}��f�ؾF,�g�g��9jdsV�1�d}<Q�^l��67�.�Ԡѡ��f"��T"��I����L�@��L�}8g�%#��4F%�%wn�y����u���Gf&>Fj����x���v��AGR�����;�)f)��4�V�e��:�
�r����e/p�����[Z3��wd�,)�b�ܺ�=��>��%���)V�U���Im0{mMkL��f�vr|4��e���D��:t�^��r���+�m�"���5I%���F����~�a�g��^�+�J�_�ܼ~���9��d�2��[m�:H1��{��J���<#�
�0)]��@j)��(�]��!5�Ʈi�e�D�C��摒!"�[Cx��~�]n}/A־"O�𽂥�����cր-lu%O�u:k�������J��S�(��K����� �+<�F���֭�|���9���k0"��6����*�x�0���4�;L�R��RU��q2�̶�i=P�L|ѩ.UxXU?�e�
6M/�ofz�7&�C�����eA�q� @׶⚰v��$<�`�C�N3!��	�,%�mY3�AF�,W�=�s@��ĩ�w���dŠ��5�;�����38/�։Ձx-Qn�?�bא���b�C�O�H���@W9-\������\e��y߸�4����q6��:�Fޜ@P�wB!��z> bc/������ܿ�6	r�l�+<i��=H ��+:�k:b����Ƨ�J�MTG�ټ�[�16{�y}Yv��"�v�k�&�ĉ�~iG&Oʱ���Y�G�k-E��^����� C�.��n��k�$�^ގ�-qu�|E��HV�N���t��;��
�!�b�@��z�ٮ�l\�U��"Cp����/��k��$>ʐX���(�܆�s�7�C��R�	��|��h6�ST��6��I�a�a��=}@PB"/4њ���،@����h6�b��ԩ���&u�^E��<�����J&� E �L5z��d)���1y��v�Z8����5\��%�}��?��w�w�(�Y�^�<~;a95Hޝ�5�4k�\�Ç���.Y��Y��3��7�g���
��h����|	ӑJе��X��n,�eO��� Ի�-�q���[�*aVE#�^�<L��H�N�++-��ʆ	�M]x!7�u=��m]#57��P�w�wJ�2�yZzHc&�ψݣ�K�ݗ�p� #�hǟ��c�&Q&0��ޮ�L�$��Vr�F~J'��h��S�P2o�@c.�p.1�(����隷����e����H:�^�������*��F�j7ښJl��+��[F;O	��I|��`�Do��IE�޴(�pU��\�KE�B3�L�-��22��E��;L�w�O����$G�o�~8O�b�j0m�q���\Q��`ǜ��ߴ�t=,R�y�m�5��4F�.�1K�E��N�`�����T��+��_�jR�맹�@|4
CJ3������&�aDm�Cv+���
�WoE�W���6�7�ܤ��5b�->&г���;�ԝf���,���Oݥ��rwX8��S	�`��^�?"~�*��Ğ�>���,(F��h��������[.�]7����t�݈���o1���j���S�G���Y��ָH���j��U��)	�9�Q�B��~� ���R7(�-�u=*�|�o�J�
��һ���A9A���ôK�X]���ؑN�(��W��^�'ğ��Cu��`}�Ǹ�oLJ���C��k0\w@׸[{7�a�6%��: l��lb��v5�DTS�4�F�s���
��~R����b�����swf�e��2C9�T�N������zo�Џ!�T_���-T�JU;�ej:�����\:�!qx����Pl1��<PtyfL�y��v2z�`ϊA��ǒ��1��Q&�w�
D� sxId�<=U-/�A������H6�	��|�dT���4���kHZE�)�?;� l����3�[��i���T���wP`kF��Jp�l'.���J2R���֥�e��N��'Ez̻���d�K1AFB#$�,�I �i�ǉ��
?��7R�f�K�+Й�1�v�s�y!�qg��/�BC7d��p�~.yg���]I&�߬����Aq>T�K�1��/g����k��YS儶��j�nm��z��[Z����۴����E9��tK&P.��0m����
���?k&+���3#��'�A�w�ʒ4�O��9t���J��9T��,����0��Z_m��%'>���x�*��&2��A"�6��mUNH>�4���� ��[�F��e�o�}�X��S*�q'K*$�xz��oPp��Iۙ���U�k�Mde'=p���.��%����8�dqt�ݮ07)<��9z3G:(�ǧRk�O���Ƈ�|g�y�؞*�"�~�
!7F�${������É�3�~*W
[���!�#�!T;�i�7K���î�
A�.1ְIi!��y��ʾcˢ���;�����=J��w�{c%o�����-C��w�a��L	���!�V2�
���=ʚ����DT���6���D��ܿc���kI�� 4�|�g��;A�Rf��F�S�%5��_g��#��n	��Oד��V�p��h�`{�9�NeZbD�9��ׄ~��؝kW�̩u3L.��I�Siy�Y�g)oi�*�RxW��ŃL�byTު�
i�.�8���U|��b�{	��sݰ��xN�1�>��q!O�'��]��$x�0*�3�ژa/�ŷ3»�àe�vM]{��kkF���PZ��Jm�(�vW" +����B���m�
crhaycn�o��m;a���$��8j.���3/�"@l{�o��q��&�olZ�6�Z[�܍�][ ��%�5���]�/b�}� �����cъK=Jo��Rh(}�DP�����
�[ј���.�k�eZ�ПyeHV~�=iv<x��a������~�lCΗ�a�n�s%|t	+���׹9����n�.��j���c�I���b����9��]����L%ӳ���Ε���R!�h+��!�����E0��>�Z����Xv]��(@�_Yp�j�T	GBM��TT�[O��ym0炭�"{�si��	˦x�����uۇ�u�]�܇���Q��QPp|f�W��]z-2��x9�&��ϩq�n-H���<c|װ�u�GPEn����~4,t4F(���Q�{��g�3qq�-f�f�24Ed��9'��B67!^1mi��P%B�U�.,bc�0&���>,4�L�v�;u%�>��2
�lF��7՘�VXzA��1v[ļM9RznhB��TE>d,:��.����X	o]0�������~�a3����k#?^R��>�5��?��;c������r2k���g��d�!����;�
���.�n��c�|#@	IИ�¤�n��PL�»gͭ�mg2�<�4�m%
��?3\+Q8�9� �O]�������L���嚡��G@�
��<�L48͈�V���HRi�=���f�j��)�A�H� N�.8s9�44V0��dɝ��u Ԗ���Vjf���-�~�r��hw���Fh�ǧ�p)�(sk*��
jj#����gh1K�k���f�S��0T���Gi[q��F�
������^Z��F�3��L$3���!�!J����P���J�� ߛ�,j���e1U����s���k>�˂���y�G�T�Z�|���;Y1����
��]�f?B�ጳ�u�-wb0l���=ēbPc�����{EQ�w` �I#w�����Cin�E�����)17R�=F�cr�/�E�������g;�I�������JK���P;���'�}�'ŧ��Kw1�j��X�t��nT=Co��������|�B�o���!og�_��}���y�C�f�Œla�9{��㨱�b
Ӛ�4��<���d������cF�����[=Lr|�}���;�,R&�`W�Ψ��wD��S�w�s�m�ģ��P�#2��aR�^a_f]ͱ�t�n@���W��i����fK��1�9\%������ ��J�� �R��4r�I�����%܂Ԥ��+�a��J��q��*;I���[��W��@ �7[�`#������Oc��\�؅f<�!r�>"�ܦ,(��;��x��B^dϮW;�qB���8z��H�С�B;�?��@������:JmQ�%(`�S�����Φ���7�a����-�B��H@�HÅ펨���^�v����X���QT��{�;w�{ z���T;ɏG!�~2��hX��Ո`�D?,�T�Ə(?2�ۘ��|�HE��މ����|̱�B�.S�q�&�2�������Ѕ���e�׵
�T�%�@�0慮�/ޱ���(�p��Q_�B�>�\�>��$W�Jd��J�.K��7�CHu�zF�5�L(�*�����ܥ$�\�cҽjz��o���K-�������<�(j��P�m�:��c�wZf͞gP=a<�f��&���h�)�X��-�e���;�|}���Z��E-�yq�=A_����<�E�_�ǩu��LL�Gaa��v�c��00M3k�A�xZď����D�9��^xcX�������!?��ℓ`�Ee�P�~�	���_�.�)�|2F���߯�z| HI1�nK-��q1��;�i�����B�ݯԲF'j^�-��Cך-�?� /��x�ZL��$�&H\��^轊���$!�?�c͔
�Y���hj�T/�����r�w,s_�`ݟ� ���+��|�h3W$O�t�����΂�ڡ��U�oY�W��XlxVHYEB    6184     f80����� ��1���"��8{5?� 8��%�X�Gq�]bvR���m��2�p!�L��v �H�ఽ�{u�[ĉ�N8��޹��I���;O��e�!�c�e�2����ƝZc����e���_��'�fH:�/+&ne�O�>dbp���� ja6����F��n��Td�F�'�J�c���m�"� a�e��I�a��������p7�a+��G�6�Ex�7��i�$�rJ��CGz\�w��ӊdD����� �z&*jk��G������)�m1톕��Б���d?-w�+��dG�D'fU�Q%�����T�Ҷ����Į�azL�|���VL!m�bib���f3"6�c�ȑ��{��	�Kkl���� ��X�[G�,�~=�je��ҝ�8�n��Q-���jm>��Oy'��"���<����K�11�_b���z��/�nz�[ނ;wGG2��[jvY c����q��fG�]��j���e���g�s ŀt��]���H���L"n��k^$��ޤd~�p�Я�$Y�]4�--GC�,�,ԟ�E���l�\mv$D�]u��b*3\lEތ���iK�X���0z3?
"�z���)R�#�5�v�Q���M+X�1|�!ԝ�|�YS�Yq9�[�@�	NG(B���<ƀl��%a/� JsQR�~{�rڍ;�Eh''� ���Be�lq�������SIte@<C�Оy��7�η�A��?r��r]a��l_92���֛*|�#;i�v}�s30�h�.X�����~;3��dЈ�H���Og�p�Q�  Z�Ɋ	X����X��@![c��A=����)�Z@��5Ǳ45�k��3�0���"��S�#](b���םcI��n�ٙ�epZ����u��Sѡ`�b�u<��_��`�Z�Ҡ9YP&��h�R�ZV?��<��;u-�[@��X/�A.ٺ�� 

����?�ɑt��dp�yzfw,P�N�-�PE~
�m��S��=�����{z )ϰ6r���Zg�fp@�� ���w���l9,/u�T�Dd�dwvhDJ��05
n[����b=���bj�㽍��W��|����[��6}�W� px�q,`2 ��G䐵�$S 1�0�F=U�N. �E8q����:u���
�ڜM��4����oV�8�I^�q����ȈY)���!W��&0�F�d��U?ϊ����Z����"ٓ?��P��F��U0�wY�H��M���ŋ���^���?1�w�Ëq��#Im:ʹ�f�R�^�"�,:R��@]��������~���4z|�������6WX�+~Ћp����S<��	�6a=?�"��|��Պ�������a�p�����d�Fta�G��[�JJ��E���N���Y��3#����>�S.J�n���c�fL��;���vRv��	��3�I�U�Sq�>��V��0V膟:^�Z\+��O���f�,���[[�>W�G|�ZO�x����[X�v,��e`��y� �G�੬;�T��H"U�[���F���Ӳ�4m�CfGA c|b�ƽ�J�ws����cH�n�/X	����<��������cR��U�LJ�%�{<�y��{�J�A����[�-yS[\�d�p�&�s��&��^�����<����{a�·N����D+�Q��_����B��{=�!�(��ת&	}�}_T�z�!��H�.��X@�|ft���߶$�s:��ljzD�X�o{�đ��Tˈ(^;[���*v���k�N�>)�l��?~rЪ9k�ey�V�O/R �p꺮@��C6AMC�U]���n� �u���F��A�^r� ��R�ӯ`𩾭��e<�M%��5�p�/"M����!�"��0F�I�@udԏb��u�8"Q�
ž��TC�'Lke��6 qy�6�Y*,<����LAJv|sg���n�BÛ��%�{�QMZt@���r��g����H%����^]5�I��%,<�����>����ʸ��T�Т<� ���KqW��U�\�e�ο	+ÆpV�������i�������Pբ;8{N�Y�֛BKd��آ�5Kg�n���pR����sQ¬��)-�"�@�Vg�ò�:/�w{�8-������#@�M�fƋ��wAt�'��^b)����9�y/�ְ��O$m|T��:���s��O�\�g�� �Q�{��?w���#~K{l6S� B.o1�V���47�#�����G�e'��Y� � Z|��ۗZ�ڰ$����3i}u��s�֔����ـ
�k����I�V�}�[s#�Ӛ�mʻ��Q�r�>���ܪ�P��,����ȮasV�	� �թ���!�ʢ4Μ���f��<��m�i��º�4�('�/�v�b��#jO�d�j�mҒ�l^�k�����]��^�p���@_/������u�}zK��<�[㘍�逊q���d�����Y�آ� ���\�M�`�F�V�X���&N]{vc��a�gf�c�q?n$r���DZ���i��45׵|��������} ��E8��9����(���Srط��K�Ont�b�x��y��L��3�w�ڭπUÑ/(a�'�"�W�M}���Ī�1fӊ���ON����)�8B�KP�zR�ݡ�㢆I�V@�ڣ��|pXB�!�������v���5�"��)9�>���?�2y�}M�����1<C�lx� f.>�u�ͰhQ�G|�$��������c��UN~���l��-��V�#r���g���Tfl���)�T�BO[,����7�k\�g�q���u�ۢ'��h�o_u�:�x�G����9��5(�đ�;�<+��M���sZ�ͳx����!�����i��9N���x�X`y<�p���r�<���Έ���d)�x�IU?�6�������.lw�3o3�%c�(O�K�.��H�y��0+�p��Ps���}��N�}n����[����~��ο�O?i��_S4��̵������a!�Hξ��ј($��&pt_�������)�6v����5�;���;� D�iJv ��;^֋Mi��M���㐹��dN�k���sE}�l��9:\ཏ�)�����X?�*�y��͚/��YK�T�	��c�I���#g"E�z�����t�(}D�ڰ�O��c�p�a
Bg�U���K��2�Xs�0�2����UˊqƋ�kn���J��P�Zp�	�	�S% �8NJ>2��hA;�� %��o�d�F��¥���S�|�O|�N�0���c(�d��P�!(\�<	�
O9����p�T_��i5~÷H(l'�N��6��B�܌SG/���J��C�m�2Z�	�E81&M�-t�,�kʖ�XxO��K�M�R[��r� |Ȧ
��r�H���j�Zw��x���G'LƗ�X0�}��)̵�O(�>����@���Uw��0�UrP[ȧgŐ4ӊ.5@�q���-k�r��}e�Y��Έ�[�eՆ2'}JKK�M^d|f��_]=�wA�Ĝ�ƒ���Rץ`G�Ƽ��t�Bc���[�6xn�`��p�P5�d��N=q�3Hw �W u���SM���F�tm"�]74�8�+,h��׹*��F�<6T���A�ȣ���I/T*���FK}�ĵK�����D�	.������^�6�ֱ�&HX��ݿ��H��i��P���5����᪗|���SA�e���8������bE$�.\w ������9���:ʡ��c���_�R�YH��L6h�hY9��N�m[>]:�P5������k�-�C6�tS������c��u�u�z}g*ƌrc��Ŏ�+T�;x��◬��"ijɞ���~�՘���q�/Ey�a