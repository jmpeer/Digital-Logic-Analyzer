XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����k<�WB�̣�{�A����l�o ��Å镤L��n��ٹ���EU�^�=����P!�|��f?�?Qιg~p1�`����e��T*�t>)T�i���k�UG��@�pR�rOR1	��ي���<���K��p/L����N��w�,��:�7��y��4"�xy�Q���ކ[X��ū ��[�H(Ns[�4�[ ���y�w�1����Ɏ�"�r�������E^1 /]��B�lɆ�6��Pg���f�Ԫ9#q�j�*3��#�8aЃ0wK�S����=�/�_m q��O���N�3~m��͢���x���9�k��eb	�v�J̤K��MCa?W�
�Q=��1�'lT9���%��m�T-�p���M������W(���xb5C� �����eD�����t��;����d�Ң�c��E}j�Ym^SeO| I|˅����b@��%�1
���e$,R�WE\�%�ܡk���3�H����Pp�fAf�f�g!t"��1����A��Y��W{[��T�H樬pg8e��߅�����}O���������9�\<�3�$0*����<��H8i���6]����]����U{�����	t����-`�
����]*u�fÊP��e�h����_NJ��0�ep�8^�:7㮚z��B���U��c~M�)��$g�t�-�+5��t]yt�*;hIZ�LƝ��C�fN�sR����=D�y 6XOL^F��9�)IBtD�	F�h�M:���XlxVHYEB    fa00    2470��s�7Ő�)�Z�ι���;K�%jnX��m���&v�Dկ�d�P�I!s)i���>���
�4�g ߵ�9���!A��H��!��3_�n(�������uU�����/U�����nϔY�i8�嵏��ۨ�()��hnخȅ�Of˄�ZPW����@��M�:${_�*N��omd�#���v�*]��2�˛iӦ^��yȐ��h�:�L�4Či���k9K+��Μ�qws����wO�n(H:H(��!��T���Ζlԧ.b;��bA%ǽL�"n��\[u��M�71�#,���S}�,.�qw��pk
�ͥȑ��<V�X��˞`VF�>�tF��
�Vn��q��5�fMu��&\b��ҌL^bX�, b���֛�ji��&�Dд���!"�o�	3��o�'�{q�N��ؘ�+�sV�!��c�o.�y�n]*v�\͋��r����2�f���4&DYYD�ʅo����.	��(d�����_�a�!V�"��){g��#���BYoF��X&"��>��1Yw]��;g�z0�[�?I$a[�+��Y��_�B;h��Z
><F/<�?G*Ϳx-O?��L�
,'2�k�.�e�Rm�9u���}�!0�&Byu��L���l�;3�lO��@2j��^e��ر�xbxfKe��OK���99�m'�BV�W����G
&d@�O����dِ2F��=�Y��>������ӎ�\��P8J�Rg=�g"�wN�D�SL�yzc�i���S�)��i�&Cҕ�"��@��O��ul�%�B��﫚��꯿�����4�m����G�9\
�8��3��_�������������~R��U�
��嗌x6^�������F�i��	vo��|�� �5=���-=������Z��*��0����*��k�g�ﻣ����Dc>�2�/�	MvMg���Շa����ZX^5B����w6��N"ؑ���VAԳ�������#��k�u�a��^ ��i�I�}���֧g�/~�>G�֗.��@�?�'#��m�O����<8����L�9�|>)�2q�C:n����4*����I��(>ʝ���������h	0{,8#z ����$}�f/1�v'|P�t8Y��kq��z�`a]��K��R{�.T�R�yXZ�"ؕ*"k&Lxq怿� ���&z��8T�`i�+\`����;A�1��#���cB��ב���/UA]�1ܮ�~觟�ʣ�%׊�K�%�-\��J�wԲt����S ��?X�=��"����?�� �-��D[`��	��*��?Ý5�g̜kP����bs�}�"~�y���8���l3��)�p�qf���Iyk�9E�O"Ad�h�!Eo����@�g��C[^�ңk�4�&��a��f�ExH���灩���j�U,������ʏ�V��>�@ ��ڳ˄��΁�U>�7�j��jߋS��V.��
�8�j��P^w������KT�Z6� ���MW����|��W�LCH@ك���e���ir��֟��8#���Y��?M��XN%��)�o�vyЦZG���
��D��" ��E�h@�2�V�l_�[�o�P�g��	��/�.ri�y� vC�(�����os�F�.��4�R@'=�G�
�v�|cis6P�W�~��s����b[4�11ٻ�X2e�'�č ")��C�^�������ږe�sC�Ă���6蟞k���еWN>{�\|Nhx �q�n}%��D��!�X��z�k�l(�y�ߠ�"��/ڞ�_dL�����&=�y�
�d�Y�z#�Mb��E��vL��/�2]�ݠɇh��Me0Qf����V��e���UQS\*ezg~���Ǣ�>)��@��d"�{n����#&�=�o��
��:'=jR�RA3���G_<�Ԏ5:���W�9�Ī�9yOa�)��b&p�h�p��yA�ϯp|��7�Ƕg��s�ݣ&h>�E�$������s�p���p���OC����@|"#*=��
��O�b&P�h�;�	i�33�C����;�J�<vf�M�dRN�g��'0�=�R��,h�K C��,�s/\�&���0թ�e@ Ţ� ����eT}��`��9O뤦z��^Lp�&TZ/��bgo"^�ld��r��l�O�(�"a�9����˺�%����ki��r�vϵp ��h וe����$1�H9ɞt��P3Om*S�F��
D�� HC�,��T�-�0W��@�n�|e�L��J�Ph6����Ek�NoAT��55I^��$~3Ϛ�Ⱥ=�ۈ�5re-,�"���Po�ؔח�:���> ���C˶��GFTW+X�����w������49��=���K;�R_4�����~�P���!�:��'��ܬ���UI�P�����O�[Y3��obso���'#Y���x�<��"�����[�౨�A�73�*ƿq���^0dY���'7m1pg6�ǺKĸw�ix�]�o��:�IV���	����-w���݀���P���b�3f�yX$�%�5):�q�XY�b�@^\[ד�BV\0~eKec9>pA�E���n
�{v{zM9�݉5�;��Q�B����5-	�}��%i�q'[�t%����"�������ƙ^���&h�#�=x�������Z���f؈��(J�G�%t�k��
 �#��+,{O��r�� �m4��Km)��z�T��ᱺb�
�jxz(��y�㊞�{�����CЊ�"��,AX���'gV�M�{�c���Gk���d�q~��6��Q|�Z���~�H�,bq�"�N�"÷c4SC2ġhZ�"g9���x	�ba�x�E�EX��V���O�#�x���/�E�j��!T�I���R�G8o�F76Vڀm^�U���h!{�������W��7ݻ-2|YῈ��k��FT
�5 6�a��ŵ$�*���I}�8!� �]K<q�6�U����0��yTz;��.�x��Z�4��D?��?���Y�'obޜX���t��Ȇ�|�<�s�W�����9FlJлk��&"�Qh��ڍ)����$�{����9��Q��3�;��z��.ԣA�O�(;~z�)�Ϟ1PD�e���UqXn��o �ϣ�	�F#X.�A�~������'�Q��\s��U�4�1��.�=�@������ba��������6Z�N���>#t!}4�=M�MFXB�O����κX�C[{{��p�� sTt�8�v�8p&k��h�C�����l^:az�$��`̈��S �Ǘ�/�����šzDJ�y�t�^��Z�/���2��*���%���"�qhȄSt1Ѕ[9��\5�˥�[�*xmS\:(2�ti��p 	knNaJ��p��F���g������5��y���e"���8�s��c�[9m��������e9jc'���d_��6%Q�Wg��d;K�|<<�^�-��D��{����I��]�����hgB�u߫W>�Q9#'Ղ(��O�������[T���_C���;Q��xs��hs6u9&5x���o5]�F�-����I�ҿ��Ӿ��ob��b����>��c�8J�uQ���P�}��&�Y�V��Y]�G���}ߟ���J�l/?C������@e����ڷ���"��(e������q�4&��@��v���QB���7�P�RL�q����,�fD�g�g,�9��nz�[@�d'��ߜ�����{em/�J��T}U��! �nh��N�@S~WY,��-����,V�#��Ħ9o3O��@�w�K��3�WSzC�l�C��ϥb�a5j�8�s�ry��_3�ד�?��ੋO���@lm�H�Gs�p2Y��E��rl�cͦ}��*�s��t���]a7`�6"�ܛX"\\P(V�t�<�]C����msӰ+�I�lm
j,x0�3�fG(B|Z���v���봓�Dm|�U��~}���Xl;���Cu��o�._@�`���'~�Ǡ�`!uh"~P��6�r��sD���fyV��K�@QO���zꙨ� ��f�a���YE�i�d����Z:~2��?���hlĨ,��^�;��C�[֣�J3�`��L�uV��x	K�(f$�m��>�;^���3Xk�L [�˨����+��wZ��� �#��|!^{��%�gz�>_��=7�hnD�xf\&U��3w类'a��*��Em������!�I�\e�G�w�`X%��ܙ��58X��Pأ��C��s��شt��J�_�V�5�V/�:���c��UL���]��H�����<@��|����N�š`�@�;�t�t%�o�{p:����\*�ҧ����o�!b#�����b�k�ʀ�b��]
�0|&5��z���� hmm��!�S�Kɠ(����E�����O�f��*(��8�W�ժ ȬsRb�q>�!̘�6��q!s=i���X�=�4��V�r_�S�i��جg׶R�c��%t�D)��Wl"������$ŵ�.�@ѥ)�}	�y��̿Ϧ|C>q�o���Һ�خ��_^���[��#h���6"٥1�N�ͱ���C�Y^��	��@g��E8P�X�O���N'������fM��K�K�&��
ܡt8��
���d���>��z�fnD>��-���ࡌ�������T���ei��)2��n�����y��e~ڡ_�Ls��3+��(q�k{�^�=`�	�Y��&�z��A��BO�	�w�TB�83����cI�)D�S{����;c�D��[6�<��i�0����~�|y]�|W1t���P�6��c��G� �����@]���b ��=7���n��l������p%�wO��1@!��q-�\D���� _�o��*�_ei���u�*aL���Z��ќ��������2�D���Xă=�{_�J���,�	s[�"�շ7�q'tn�R/0�D�Xn��N�����Tx��/zhLD��$e��͚[檜.WN�Bj�N��x,��¥�w_̢[����F��׀.��1����:�l����lf7Jʝ��}��t̤�f5)��)�=����u�#f� �z�9Ul7*�ݯ�L�>e������5W�}J�苖�Lt���zoX1=�}��%h �� � K߉û��8�_p0��q�_/)62�WQ.{�,�"���j��.�������,�t[`�����;�I/���}��T�,ls��0�QW�>�+���yI�(��L�G��"I��O^E_�l���B��v�q�VBV]��Є,�1�͟řL���rM����:C����)�(��.e8�0)8����Y������� �y")d^㜀S��νM䇞�pF��������ڱLyY�TB���n��s]kﳱn -�Fq��AE����@��D8�g���r�H.:�?gX�%
}����lPKJ10���Eb@Xj��HT�{7�.����v�&wH���&"��!���������O�JGv�ǌ�'vS-¶?.�c4�'�!�lv-]�aS� �`
4��/���|7
S}�T����y?��:�P�I�
�N���W���-�ܨNa�2��9�;$��ξQLP��=�{3�ω�H��^�w����?�N�ܾ��ׯy���(�~�+�c,�3dBZ�݈F���z.�N����`_�@F�o��L��DJƊv>�q�\s���C����c�s��_|��##&٬�ᗨ�N&�F�bB��������0f��	M�T}t�iW�c�ȊU��?W�ƶ��=kM�@�>B(���n2~��!~������_�YL��բg(�h'K�GouBH����ư�=cM�b�r~_;*(gO����.M۹���J�&*a�+{<�6"�tH��`���D$iW������C�*h-�ጏZ�����%CG���g~��c���r��\�[#uTo������{ު��:�y�O��q"�X��n�ve��]��=]�Gc?��w�%@c�;�zO�P�Td��)"n-4��*�Ww��g��e��zPh\�$+li�a����b��x��8�W]�bbZ�=ͬB�����Q�u�~��7�	S�m�H�߃�4
���Y��aA���(�f���V��KKg˖�if�H��2M*5��������ѓ5�0�3M�b�G=+(xΑ�t˞6�'56��%��߼�TE��'��ea��4ȹ�!��O��L� ��ɔ09���v��TX�~�a�����S�C�uq\�t����I%�*%z\T���^��c^�N��������ui��ʔsT�NL�瓬S�"'��mt%P4l�2��jL�V3p�.��A�g�����W�
,Ju��M[em����l�� 
��#-�;|������N��!)ї����`�z���?�ZZ{��l(6���&�U����Eh���9YE1T�CHꕝ��H����S�T�3R��Nh'�T�k�dŌ�耶�RF��b�rq�#��a�'�7�َ֑��: �1U�Kj��+2�>� g�1�}>�ҳlR�pq?&��	�(I����H�[_.�mt�}�+�T��W^���Ձ��ut?lc��o��>x&Z[
�j|VA��i �"�٣$0Bk�F��8+�����[���[.�#ك���B��!N���h�vt�a؈�]�,Ӎ�a�`m]�Y��� �&�p�l]�$e=!qp�{{�|`��,��f�;FR�?^�n�{�Ξ�]�%�+��Ԓ��P_i<	+���P	}�|�9��<,���U�E3,v�Ϩ���_M�]�=���+k{qiADb�
wɞ3+J diay��PLr&��&��"��a��9�"o�qX��♉�����n,��<W�.�"�
Ԙ�@�N�fg<f�!C�[3��I�� /�"vq�7��ń����?/�z*x���l�������j+N��{=�H:�̓��2V�5�8�ѱs���'~"�|��v�	a��l�=���<?��S���F+��b��yT���]�� l��Ś��*�t|�������n�*ĝ��J:���0��oq #�>`!kI\4թ+D�k�l���*���GJV,q^���=9@-��8T%#a�C�X/�va�����F�
a�%H�*��A>�/L�v���}�1�<#���S����ލ�yQ�����1�$�7^Y�
���)��GAv�@���2c�ko]_��Z� ¹�H��(�z���f������:���(���;Gq�z�[���1}����=3�$�a�V��3�1׺��{�_I�
���p�~'��۶2��AK��1:����Kʣb������q#~�!���Qp ��=�#��H� zC/�V+ '$���ծ�dêÌt�̜� �}M�;��Z�K�^0��"Γxc�������{��x�8�:V����y�;ή�-�����6�( �+��UI�f���?��X/&1
�Ô|� ���6�Bjo@�Z�U�&]8�8�1�4��󄵒^�P:F��k�a�+n�;��̒��PL�@��5V`�Њ %��~�N59�5٘�Gu�e�-��>܃�&	��c} �����'�h��V��$��k�9+��s��]�Y��,P����⋼�Ӑ4�-��ݱ�;0�61sa��,j�����ܛ��\ⶔ�X=�=�#��="��6�uf���r;˱tom����:Qdı�E�t^�w�{���~<���ki,t���\Ϭmu72�oX����X龷���+I���j��F+��t.`(l�	�3
�pӋM�)���(�ϒ�J�-%I[|{�I�W�F�݉[��(���!'R޲��G���9#SR�˴S7x�/
����\t]�le?�4m���OJ[i�و�#$�ȸN/�B҇�i��Q�ύ����H�:�?o2��ߘ��j�+繻N�e�UsAط�Hq��O]`/��!�b������.��{R]d�U����%r�Z{���E��\*Y�&Ty�X�@���>�Rs�P��k�z�ӈ0�A��N��P��h��]{�.TA`	�,:�!�+����V���)�7��,8��� �|-)�5��ܛ}�b���%΀$QE�T������0ט�<�u
�\hC�4g��v���� k-pX�eo��zG�$r�Ξ$T[�@�
}�":�����Kj0�����W����|h�t��|$�Zs��B{�ɩ��9ࡦ���4�3X�<���h�GQ�2������/��z�����8x����[rC }e����Z�[Ƒ���9�V�5�cxD4�4,@j�:,��
������e9"y6��j�	]Q�;�88�w����j��c���f�wi��ig�9Gn�~ޛ�}F>�����`��n����䯵���0����Edؠ/ޙZF��=+$��#� xd��\�7z_�[	v�x+{�D�S�K;��a�LV�H�	��z�σ!bْ\I`V���z����e�H` j�"�A��3ݰ9��}�*M�~�:�Íz�) 6�Ǵƴ�s>�p��	� ��A/Ѵ{�/���5�=�Z�i7��'�8=5e��J')�e��^���z�����iN��,P�а2��D�`�4�v����0-�U�kf��ƭ�X ��y�#���D���V�U�Wa��EQ�����x`�E^\ٴ�:�[C1`�P�ȅEӂ��@nNh�f��BDWN��r¾,H1�=tf�qwkk�\3�Ю-˃ERl����v��F����p�r�n��{��v��KR��n���b����7�w��X�b$�3 �Z�n�<�g{c?�����)�=�� 6��p��!P���7C�_��gT�B��RV�� �� c�5�+�ў�Yg�]�E7&��O[����t�ik��T8f��H�&}C��=y��֎8"��#��,�³�z;l�6g��N�y�����Rs�\ؖ�0��h~��C����Bz2�c~y'k��:��[�G�?�pl�4��(J�����(M� �B#��� po0f$��Oy�i�\^�٤�״�T��B��/sf�7�����\����_!x�N7:w���G��Y�����1G�'y��c�{����V�Ѐ�7�ٔ3�%�V��y@m���Jg�F�s_��[2���XlxVHYEB    fa00    1b30A�=�glR�u�}����_��"}�>w�3,�V�Q'���c���ko	B�F<�9��j>�&9���X�(?#��G_U�Pϛ���=�x��y�����P��FW'���8�p_�	t�sn'���DLqA�\=czԲb��!zI��ж�w����������gY6�7~��9�*����۫6��DX3����n�y�mS{|����BA1}�=���>�#���!����~1���xt��Nz.�q�X�3�~$�`S8�ԝ2���A� Ҏ|w��UB�p�G�ԼQ!5�}L��3��Ĕ�2Aű�WRI���oF�Թ�gYտ�*G�c(m�v�! �j<��`�D11\\.E��3>Ǧ�En��S�U��7����vB�@؛�89��',���������El��+�cM�-�����G.��;�}�#��+$,�v�ہ,��"p$e�Y;��S&(�Q_�U!���t5�yŉ%(��E�=�n�����A"��wIdZ�|�?�������O`t�eꄄE��'��U[��Pǅ�n�y�<���nJ<���?!��s[�εVD��V+�(j7��ufj��G�B�^>�;-)���tb�����H9p�rj V<T°����ւw����}qBFb��%����KWc$4��c6a�*���"`���F�Z��E�/��Hj����79�O>��`�� �!�5_zŰ``�#�9�Vvi�ܛ̬w�A����8�%5^���az\I��8����_?���.�A�4��)&3�6M술���|��I�Zնg���e
}3ف�<��w9T�W�C:V�"O�z,�"�v�\(�B�Y�VZ4�-9�ɮ�T��w�Ͳ��f��*�K��v�:��DL��	Q0H$v��/j�gM1�O�wp$-_�R_^�k�ޯ��7��fM�(�iZL�\,�,e�iA�"]C���J`԰�i�f�����o���E"���Zgc?�~D�:�*d���^��
\١EM�p��p"���9�}�o�i���pR�y�Α}|S�9��!W��y�3}�]�²ނE-
+qG��*�����!DT<�I'�]�
	۷P��d8_B
8��A.� �ɷm��񞰼���������G��c�{wKO��ݖ;�F����C��V0��̏7ξ�$����$�Y��6�=�OWt٘�CY_.5=|-�ΔeW�)�&��ݰ_�\}��H��^�.��8�O��,7��'c��y:� �s���$�&(T����J�01����Y/�y?�e���^;�M�˔g;���ĝ?��`3*X�Gk����pz����O��"0�۟�C��ݷ�<;r�u�|����3Xٖ�J�^-���d�Z?kH�z��mH�V��_d�H�=p!`cJ[�����'�˵!�k_r��V�2=�3e�G��>�\��f�i��G@�H��S\�s��*�e���4��&A��Ոl�+ƌ�T��=z݊]��t 4�� �:���f����4@��|��J�M��;�����je����;�ګ$�1Fm0�e�����щ��BcA�7h����>.�;Z�A�F�_�׳ ��d��n�tq:9�-nLᓛGSNh�Cz@�/�7��Bc{4��g�����B���@7 <������=�r�p�X�W���q��7J烡8ngv�1Y�z�?�ziU2��,��@��� B[P���X���d.�Z�״l���K>�<�����B��e��|R1�kl��Nv���;�l��o�{d�ف�����TK��np@.ş�U@ ����P�!r�j9��Ϸ������l���~����7�� i�*�x��v���j�y�|���V�`��aлw&nc�T=��Q����j=D��4��L�X����yD�g\6�+�W'�ؖZ��x<�X����P���[4�1�`+��Q�?\	�@�H�̗ȷ.βi٘���eh3������]���g�]+X������P�?�b2��yy�px�Ȭ��y磕R1�p�鐶�_p�[��p_S�8Bѫ������<�t�1���C�޲�1�u�eŕ��Nʦ�w��0���&�<,��E���Ű������5HL�G;a	�y=�̈́�H(
��CAD�����Vp9\�#��T�,��{�Xu�
�P����ώ���d�(o���[�QB
���<�P�X�ob�Wߍd�q��Bxi��8�9�qTZ��I\�}�ԩ#�^�f������P6q��Gp��Kf�X��g�g(�sz7�g�_n+q��	u�G��zQ����o���\����Q��_aڴb}��J����4GE2�p3�W�8�!`�h:z��a�v�
���Jm�)�Nx�E&b1���J��o3~���gK�[3ʼT�*x`��e�C94��I��WJ�)��`J�[�(��g?X���!��p������y��m�[~����p�Z��q�a���	W�>�ٻf���{�Sf7��"o$��^#z��%Ԟ^�v �"6���#�0�0��}q�/ #%A��"t�y�b�@��V��ԭ���ے�Z��h�%��ȼO|]F�MS|����y�ڶ�1��nl凱뵣Ҕ�r�!��+��Z4u��o��.Yo��W�E��Dr�BkҖ��@�L���U�-hҰ�?��>�uHY"��F�:|��O�5MV*��:c8"(���V.���'����yJ�H]�E@���O��G���O<x0U��_j����s����s>�?R.��-���z/�̢4�k�@J7K�G���n˘��ݓ_E�6��N��V=#��=4 �(=���D�r��l�Մ��sK��"�+V�@�Etg˄�Q�;h��+F���z�*c��mI��_n���_ȅ�,�����4c�K�)��k�^{�X��H��n�-+Y448%��h�"�9�#Mh��R�����'r�ܬ[���	6���P84��
��&r��:�^�0���O���D$�d���_�v0�=+�?����X{W�DƖ֛��"B�M'���n퉈��ϥw��L�N9��X���in�;W��'hy��W�(3�|���E�#w�����Q1fUb^����uړ�n5Y�{0)�12.)��$�1��z�����F�Vu2��i��Ipn��/�nɪ�l0T�s����4֭6�>�w� R۴Twń��d��:s����{��:P��r:+���H�G����u�b*��*>_н2汼�5�ު�K�����mO$Ό�`.&���͍]u���7H�n��Ě���)V��+��Ӕ.���	�o�!�F�)`=K_��J��c]�V��OT}^���wC�	�;���"��3��}0�{�D�)�߃�d��'aR�I��K���s��s���<N����\���f��GT������\�._^V0۾�������z;K��Ū��LC_#Ȳ}�}8F�!�kV����/y���!���-��l�2��`EF`� ��"��.�ꢭS7d;g��x�9�w�6i�&i����n[|n��`iړ� �l�mL��h@?BV��NQ����A/ܶr�� �F<ae4	��fD�<�\tΡV{(#	��V�í����)I���d|n��2�;~��m]�	��d��s1����%���}:!g�����^� ������;��R�hz��#|)� s��������O��o��H�t�	O��|��*��e�Z����C&`��ĺ�'���;���7������Fì 	���_<#���H%YK8��vdY�lrm2fFD�L�I��`�AԒ� h��?|~4ь��ma�����lR7b@n��-�~P�=�ds׏	 O��W���DV[��Aʛ�p&f]����p䁮�`c��3�0�-���fd��>�}	8�'���p���զ��q�MN�&�����`\Gj��Q����H2 d-���a�tF�|����A#��C��8��}\�,g���i�ݼ��������މt��`���ő���Xt��8s���O�g�]����Ҩ>���-����z��sK��R����`�8��Q["M�%;�`L����Wa��.�N~5g8&S�A��o<�΀T��}2�ё�}�e	^��~eǸIC�>�=oט"w����B�*7���$��k�d�dn�쭮�?^��y3�{��8v��c�������\����3.ݙ�PJ����Pv��{�7��3܌��j�����8�+��U�C�,:�10��^�����aId�E���W�������:�a8\�8y!W|q���&h�N��_�Ӕ��9B7�Ǔ���M��������A/G�@�A1�L�_���#R��;�8��@[L ��ao|��#�կ�ʋJ�R���h?}6e�HN��3vVؗb�4������̟���R}�7��!+���ԧAh��v�]Y�}5�#b5ÅCr��Mtz2ǹ�LT��%���"y㞝�$�8𽃜�k���K�90�^#���$\�d���Ŗ=�,��t^Y�D[R=d]���pw�2p��q�ı6e��ۡ�t���w��xb�1�S�<�w�q���̍N-��ÉT/��{�5E7]ʃ���Jr�?��- <����>#�1�?�IR4 ]�����;���/Xɭ�|ST�y���S�{C�'H�u��ͺ�#.��Ek�bz���ت&[GYH���o(>��0q�Y
2���EC���E(���uʨ�4}��-W�ő�"�pb�Q���q�X�[52J�P�c~�MDJ�5���&E�Aǭ2�Ŵh/�묞:�׽����O��So���t˾���ԂVLL�L=7 �v�A�(���ӻ��h~m�:��9>2��:)���"���I7Q8c��<�4xO�.��G��l@3Ʋ�&5���-R��X���y��^x��r�x�.�����V��M5�l�mV3.r��-&70M�QLL�PC�O�'/u���;�az�yE�Ҭ*�-i����Gr��bY�5��G��b����ْ�~&�-���0�����WccU�眬��-��V8��Z�,�Xm-ƹ��x0�P�T�#���_��Rd�XHA;�T�&�⧺_���7
��L�D�Zϫ��YWOʡ5>V�/�.��Νz� �B}qo۾��[�oOrM��=��=֓E��$Ԋ��1�J�a/���Y�}�y�ʂVP6����c�
+��oUed�f���FOh������p~��Ю:g�St��y;�+9@>(���&�9�SC
T·ڄ�@хj�+��)��@�ʙ�� ��/{n�L�
ܹBBO�v���m��sž�dX�ma�U�^�f�R$�.E]bh�x��G���\\ɏ�dy�ii���ژpBV�gM�]�1]6�q��/�29d��G�T�T��������i4��aC�C�;W95-:����!"�М���G�� �M��I�`k������KRٕ%q�1;R�Zn��Fq�W�+J�����+���15D���^�D��Sx�Qw���w���7Y$Y�gI�͜BP���v�>����*Ʊe�K�8z���N<0w	���`O���#��~����8�W�Z�>o����wŕ�A�'��n^������tM��7��y�M6��v]��O�Ga9
�����e���M�H���G��9�x~�m��o�L�ܯE|�2��s!��fnȝo	>'�c���ф̼�����j����{%���B˥}�TQ��]`,v�>PX@u>�V`.^�-��]l��39R<0t�8§:aR��B����1a���[��F+��2�^�5��Zr�Ƀ&��ӻV�L�J�R�x���U�c�NN��`��jT9�v��2p�l�ѩI�q��x���8a�������E��`��T�4�Hc��M8�9�拺�ȫ��mj���Q�m��h<�<Ôd`Y^�x��q�~`�M�p����'Rk����N��*p��4���W�����`(�žf�M��Ms�����6���g�cW�9���<�6З�[eo���(�)�R)�v�������s"w���/,x��&�֒����}6i4��9�EZ�q�K
m�c��pl=�t����ZRm �p�Ł��r��[	3}�
�<�N�96E��9��ճ-	lfL�$5�ۏ�n�"��q@y��qJR���ɱ�r��g��{�彝����Ε�?���ȇ?tߖ��gGvpvb#��ï��2j���հ?Q�%DZ�����\�Vk"a���J؞�*��*A�h����W� �t0�p�';�<��c�!i��0��%]�r�~�鴏�|p4n��dz&���[_�Qy�s�1�D�e�ZeW�ߟ�bmk�_$r����De3x7�4�B/��{���P)5a�j�W��j-7��N�ۛ�����5�{���â��@�Wa�M�]�R����{|�(��*����6˓x��Z������o!My;��A��ܽ�U�5�pxc�y�,�I��
�`�o�m!�_۶�ΐ��w��3����P���U8.Aڲ�U�]��Dc��x���,��6� ,pc6R�)�^�o:�kL��&4���=� ���I%���)"�?D
!��.y�j���捨f�J!~�qz:�ҕ=?��K� !�u��"��9[���i�V���8�s}̶��"�sBV$䇧�ug�P���Y;m�� 2w��� ��S�3�]�8��\����q�"�N\F;i7��,�ެ����j�6P�s%U�6!�}C޵�b�]��=�u6�z�pz����n;7����>�QW5uW�_iꂍ$R�H��� ���딷�XlxVHYEB    fa00    1950Y��s�]��[��U�	VЮ�j�Ipi����| ˉ.��9�x}����
�$��A|�o:p@�O���,^k��Z��S���q�2�𚨆���O�(�y�����`��u
��5�[����MPn�j�l{G����|={�2v��%w�?J0��0p�~��_i�^X6�Y���g�w����g{Aal�tdb~�4�P�j�fS����-l��2�|U�pep&w6�f�&O�lwdL'"��3�a��/��V�s�6%�V���Ië�v�]ڶ̈�'��	������v껊��.�͹���l���Wۿl��Jci��C�t��o	*g�KA�j�ACF3=�Q"Z�D�*����2x�>D���vy��*�/�8_�]MЁ�Yv�L'g�0gƵ���"[�	>�ct=8�� :�m������^�����}�G�0��N�܏&���!_�&6�':=*��[[�Aʆ{,&yh)�2V;`$��De��lq���bn����Ҽtȍ���'}Te֋�N����a���L����Z��Se��3��TW�5�bg��\D���qΒ_����Z-d�t���'䖜��볡-Y�<��Zy��<�p.��){b�t����1���w*��;��σ���u��w_v=�V��{614�C>o�
�Jً���`�+B��t��x��}m��W���gPE���x1��H��a�ڽ��E��B��*w���d���_����@�Q���k�D�0G>x��=)��S�e�Q�#;c½$Ϋ��ǹ%��ŀP���F�_���AI����z~>s���&@�쏱�m�� "���I�C�׭��3 ףhU�����N��Aħ��Gx� a��d�mP�����H� �eʻ�8"p4��0�c������p+�U�o!�H�����S�H��"lZ�Vߓ��27�����c7�X�'o�z2ȫ���t�dYL�M_$�T!�z1�NMC��:i�P�§���Q?�@�~�����œ0�ܺ���m�"5s�=Ţ*��p/^�ާ?s��(2������ɀ�p�C�h[�q�ݧS�� ����5��?0���-"n�od��^n�A���'H��VnM)rN������$��y�����1uϪ@�EC�A�uK��:�$�t�U?����) K9ո����&��¹{�/ʴ�Hr�L/cEH(-H��zm���?�s܋q1\\�]4���tn��C���£a��M!�F� I�?��P?;MR��|L���א���U�e؟��XO������WDU@B/�6���_���d��xE�m��ظ���/�&Ѐ*'�!JA�#��5gj%��������5ԏ��j}�㏹�;c	��Y�<����C�|Q��t�ǽ���-��:؊�������ۿ*��u�bns����"`D��N�L]�;�R�2$|Ӑ:Y�fHpv���,�>G.��m�����m��rh��[�y��1_W,ByT�m^_cCW�I�o�Ѻ����Àux������M�j���/D�'�XS��mT���T��b!��D�{Ĳ���b��:w#mUĢ��Y*ލH��Y9���]�Jnl����-�Y�`_$��98�4��I�Q�́�G���2@��m�;%Tc�~�'W���zc����'E
_*��.F?���i����m�>���u�t��S����%���j� EDNu�:%Q��*>��%�*�o��aX��a/�&of�=j�{��sso����rm�꟣���zp�����i�|��s�_�QL{��N�<L��
A��Cv����yF܌�ywY�]�:�m��&m�q�i��@V�Թ��<�W�"�q��y���d2�UCo	�M�-p3޳}�Cd'���Ev�@�<L)R��G�\�H��PW���C���x������r�c8%�R҈E�qP�@�� J��� �M�p܊Yyp�b{��;;u�vI�?����w���뱒-�5������f�Ar�����E�p���Ial>=XLߓP�3��*��G)��_��}���#V�Æ�q�������#�xe�S�8�E�f�{i\�V1��vns���K�4��,/� 3�!�ߘ��V����-&W@p8�����<4�Q�WOK$�J��/~�Z�:����N��"�[���G����bP���������ಪ2/v�@��W%�÷E��pX���k"�����$���Y<��5�*ט��ćO8Î�C�	Z%���Ǡ6r2�8C2@�;ዺ��q�S���aN� rNy�{4��,M2fp;4���o�B� "׊y��9Kz,R��2������\�#����7 ��4z��!�uٝp[�\y��ـ�9����RpY��!�:��Sv�3��|Y��r�(��*J�${θ�ɒQ�(<�Q��K;>�nK�$��nK���Mt�E�Ŭ,-�0�I�]j�T�������ܑ��ѧ<]&i�T�y�Z	�����tz�ʜ#�j�(ܡ���x��
��na���xȚ�W'9�k�b���0��Djˁ��zV�⁹_7�(HL���� �[�	�>L�����hC�����M��%�i�^���⢐8a��J����"�j��L�ܹא�R4�e�'Cy��]�ܨ�q/|�񆾏a��|2��H����r���+F'�G�[��c%�����oF@;�1Ӡ�L�R��#�PDU$�Q�.ai&�k��N����Mx�*?�e��F$��0�A�m~ �S#�;#�����0M�ҥ$�)R��^�ܨi�v�Yk���ʄCC�F�*Y%!�
O���Q]�̡3P�O���� n��Iy��85sQ�?���k���Q3Hڸ�R�b��H�i�r�R/�6��ӧ�+1X��� /@aM$�D'�c+�{	�-���N"<�{\mj���f�������� b"
��P�����M�[Z:�?8Y���sl>��TTH�ds���Ύc5��vo�])�4�����9z�wxN�wB�J� vC�7	l㋗�4k����q)����x�T:��B'���+-/�a�b���b�7J�t�L�D�@/��\M�i���svw=�;侗���Y�?�Ȯ&���!�E��K"k�ͼ,��<X�uı�[��
���@��:���U�~���@s"Wpet,��+�?��iG[�l�+�U>��u1�o�����^������4Q����,Q�����I8���j�;D����B�-b��+u�Y�"���5ܥ�3fP!a]g�W欐8�P^�CƧ����x��Rlb��!���b��q������4�'J�'4���ܶ�{F��T��l-5��ڄ"����A�L��g�m�eD�`�Δ���+�5�>jQfV��;�J�(\ˎt�t����g~ע����~�j�k /��u�|D�����&���t_|*�"~<��)���"�Ƭ�#.�+O���!E�i$mڌ3!�2b��I��"J�B��OI�kIZ\
'�:*A�Ʒq=�I�Ȓ��̡���4���T�d>5մ���ۑ}-���D�d2a�+ ė��&,#U��,h�����S̛q�;��R^�(��^����IP�/R���?3�v|��ִ�~䶀B�t���}�z����G�e����|��V�d��b�+��Xz�L�� !��9�/�u��U�E$��.�(hc\K��,ʽ�Q��<t��W�Ϋx�I��[ @��i�Zկ�OtE��e�	��YИ�n����u#��ǋ�	�}H�'���K��w��G�e��_f�bጩ�M6e����
ŏ������K�(ݘWF�?@�	#:�@��c�<�Foi@��C��*d�Z���<3�	&�/8r��C��؆4�q�ݎf����[/�Ez���c<3�5��m�Ȝ�
Ħ	�V( �6�f:��h�SΐgH*�J0��
9�R�� :����q��}��Wg#�:�
h����
�&0�w�1��S��������n�����n��:����ȃg������}9�z�Y��2��@4ĸ��4>�ϻ��I���bi���)�|�
���
:���e8��f�q��u�P1��/0d�=śv�f!���53i��//)Y�1T\$�D-h �*�@�K�[ ��(&�9s*!�O�Ĝ��^Ğ�c�v�׺v���^_ˣ�M����7���ah���ʄ�źap�_L�Zww)͑��L�z���앑J/]��yD���`�_q��x����&�8+IxE��~o��Y���u��,9#y�Xٹ�ɽՖ�����>�Q!s�E?	�V�c�K2)��O���2�����\{��&vdM�+�{9�Y���2v����f9m� �F�:$�.��	ľ$��Or�O�W8�6:��7"] V�&�����!�G"�i�ղ4��X�R$Oʡ0p��'yl�����&�p|����\Iiu�^a�H ���rm[�pM��>��"�hE�����C+0��n��<Y�
��"��3؏��v�S�����n�~�^J5OR�"�e)F/I֯.��Yl4�Ʋ���*j��t/��L�bGkaQ�r���#P�:4v������?��FbjT����//(� /L�^^�t	t���A�ʓ?������*Q���T.���F&Q�9��&G�8X�����3}���X�3<m�} �M!�lP_'�Mnq�w������k�����~il�=U=��e={��Z�q���Z�����x�Y�!��T���a���u֤\-�6'��VQT.��׮U�k�G�X�%�B�Q�~z2��S�v�7+�t���z_��&�$�K���Ƅ��a�D�(�l�u����ͯok᭨g��` �+O�0y[B��$��[�2G��e�i�U�r��C�s���}�5xM3�Ȧr3mUfaL��e�s�Yu�~��C^ Mm���PCtl(�!+�d"���&'`�U]�[��	a��Q�{���O(��mV� ����<a	��`�z��q!���f𭢂ݭ����1g���sç�n�w��N�h�d�3�3 ����趐Y31�˧�݇��Ո{����%��XL��-����g7�x]���T��=|;u���)�+����Eg�ƒ��-w��]r!,ù%�g~T�M{cF�r����~눞��l�%=I���_$#ȱ����r�C;t ���t!��?��J��.��.������>2z���e��=�kǙW��דS�q�vP���=r�{����ո�?L�+-T��8I����@U����|p�Aw�;c��h�	l'3�N��o�|%^}{|PN�g�au*x��P�X�ToU�&:�9�(��nlA�DN��ck�?����
K�v�ǣǡ��v���)Y3��/�����blǮ`�$����giy�. ��#�.V%��~]��%XR�ŦB/�7�?8̧����9�T5��FG��;��jd;6�<F4)k�󉙴5�f\)��i|;&�u���� ��Kƈ�ͪ��!�����S�z��y�ԓFN��������yt�����6/w�qH%����"drʿͯ�����z�����pWٸ�1}B��U�и<e��N�ܡ-0�A���>�A�1�|Xw �ʫ �O!�U�`&�if�����Rd�i\�I�w:�-�zUi׍=] A',t��7��y�S�H���?�,���2Ȩp�e��قp��OCl�n��k%�>O%G+��b�o�y/>د\���Ж�_+O��_3���*��!kpF4S�o6�nr�fhrNc��|J�ٞx���-ά	j�k=�Hi��pt�
M�= q�˱!q��0=�*�
�LБ�[��b8��b�{쮐Ϡ^t;�KZv��������T�H�@�UF)�A� -( �%:=�ԃY6*�F��w�����>�����'����^P\s�_��>�EL��ſ6I�ٶ�l��e�
��V`��8��p��L���l��b�? ��C�I�8[�@�J-���4�����X��<�ph�IG��԰����f#���0����բ^,�����) ���\���^�¡�hK��9�s(���������	Ҭ�i�YRћՖ�W�%T��tC�1���3(�!4�pE6K�����r���q�^�w)��u��2T�s��'h��N�E��ǱjD�'#�9dw/�7�$�`ۍO���!�x�X����9�z�.�ћ�Ug����op�"���u��ٹ�B5X#m��@ �y4���:�Y�c��H��1B�v���{<�!X�@2��� m�1�A�R��=j�����O_���S]:�*��:����m�����7���;��`���ȡ��J�Ap����M��>��{XlxVHYEB    4f27     d40�����C�Ci��s�Ҍ��Z	f�(����(��'qr��&�޴�R�@B��G�����y N��d�-�/W�n��j)����:ҳ蹆 Z_�E����(�}ԛ
�i0ma@��@8�����#.�P����Q2hb۩ʼB����586�s�vu�{�i����ʞA�3���<�C��P�S_k���Ki���9T��	-<ĳJ���@J��5�����B<j�|�O���Ԝ�("I=��Č.��B���oF���/R�*�k�zľ��$ �G �8�8\C�Ͻ��~���<�w���+�y�С!_߮�#��N�@�=gWvF����s�V��5bB���Ԏ���>m�ˈ�1�y{�|���|��N�O�L;����.���}<���~����G{����[95����B�� �&9=wO��]� p9�*,Z����U��+R�}dtN�`ƽFe΅�6�Q !���S{�o��u��ޫ�jy
P����DO�ެY����D�e���`#�%���ˎ�U?S~ï�f���*ny�u�Yz�|8��&Ę߽�Ӫ�q�^���L:m.��k�-_	6�É�_��r �(}����g�0�~����={��H����^�Gs��Tg����n
�=��0�W5[>����-ѳۊ�X�A`�^+4T�3B$�,>���apV|RH���"�kz+u$��1��אt�ӳ��J�B�W^0���3-�d���w�3C*z�h�E��KM��Z�TH�����)]�@vj����|^�'%C���!zx^&�tx%���u�t@?���n��D�%�5�/� .�n�#��	�Z�y{����麵-�C�w1���N�?^�Ęx3`����ż����X�Z��\�U{��"���͝�\)d	 t�(��}u0����t��M�Z.+�����c{����/� B�7�*�t˩�i�.*�Nxmrp8�&	�VP��6|
��`%�?��:(ѯ�l�Fs�d�����D	D�nǢ43�����j��z�U���|]蛠�\W8[�kM�b�9��ox���J�ֵ�l��Ϲ�45.KDt�Hl��m���>�������)�`���nH��.�Je^�ZmPKO]�F�{�%�= ���'nص��#?�FCJ'e��C*��^h[�-#D?p��a�����̽4�=\��a~9r���	����zXB�MM��I6`��R���T�BP?�L2�4r%���Z �ަXF�;��2x���̩�X�W_{��������Tbq�8�V�?^�>�-������rgw���M�E���zf��d�� �.�e��U�@�o�^4�x����7�%�ȅ����?F;���� ���W����@hւF,�e?"Ζ5�_���&?NTT��f��%���D<�ɣ+׹�0�G"�1�\8����6;���'V&��� �K��īڰ�`5N��~Q����ӏ	����훴P�S�A�d2��'�
K(N��n��C��@� F��t����6�X���"�<�e[@N�%qT�/��*�_3��C�����\��SO�-�t�Z ��\;�))���W_C_����ǘ�F/)�.�/v�G�67���^��Ilv]�-M�����Anf����`l��)`sɍ�G�ʕ�4���iT?cO�Wpu�K��S}K�_λ�y�gW�m�ܻ�$�8�wߢP~1;���Z�����2w馈zMʴ��5F�
f.\o�Y�2����RO�$M=y�r�Jzշ=�q!I�? ���X���Vk��K� w��5[;�r�b��S����S@��j��pq ���O�7p��{�:��ב��Ga�1��!+�!����h�hr%���Ԛ�9�{Ζ�d��QU����T�=��F�3{����x����	�"��#�3o+�T�3��_���2�A?vmb[�k����;�`�"�34o��w��q��J��x�B<��F�Gk�}�b�ݎңB3w�Q�8|�Wh	=O��������T��<(�bL@��Ǒ�9��䯤����.g�+[>�P�=��2��",18�6�1m��ǜ���B-���L7�SMG�=.j�W��&��b��$�C�{h#v�P��1��V�>�g7h	��7!��f۞�/�']�3
��_`�ǎ�EM��
�����D��`�#��xZpXg5�qO���E..��z�����Y��2!cXA��G�`�J���6��P�.c�46�w�mw�+�KF��Ȋ�_��g��� ^.��[O\�;�PKz�^?יSH�\��@主�H��������rkQ����86i";����.��ͮd�5 ����-��f�|p��	�#H�/~Wǃ����Z�{$�!����$P��������~qh�ʋ���tn�n:R�Es�����Tժ�U>7�A\��«�tRH"��R�t%���2�X��Ϙ���0��} �M���lg�o�6g��ƗJ�����;��̇5�ǲգi :�yԲx�p@�"��ی��:y�`XKS�՘�B�����u�Sw�?>}<VܚYz��8�$��f� Q@��s�_�b�x7�[#�89d���'�b�b���GE���Z�¦�?K��3�B����B� ���B�g�Hz����o	|Vo��S�ްSJ���!J@���p��jr��@��c�D�/q�s�O�Џ���ъ�?C�y�c*�?pǰI=������n�x�˄��R�)��D�Dn�����]��/����1X a�9���;��և���SJ�}�J%|�^��n�z���y iB�:{�O�t`ّ}�?�]ʓ�`���T�\�	7�)��_q�4z�
�ț,�����.h���f�grkX�K~R}��q_1�hh�8�Rs6���;(���O��0�rytJ�<�qRV�Kw<ۄ�����{�	!x�4�A�t��)�p��0��խ4�J�@C-�$^	
S�*ה�_�	��3�<4���pq�VU;���>�{�a?b�^�(���-��؊�tS������V��L
��A��g�w��GwNp��/���`�0;9ݸ��A�s+�m���éۨX��`�L��"��!��̫o��@i��Ľg�S���D-:�B��-��j ��mV-�!�J��)oILm2՟	�%�?�N	d�_�f��-�\ u����V^ǂ�W�W<i��VD�++ ����l��]�3/���f�h��R�Rpe7 �#��%[*�LW��cG������9���Y��sV�q���q��]��}?Ep�c�J	0F&-�F�%�v��������(��z��&��9�Ϸqfiq�X