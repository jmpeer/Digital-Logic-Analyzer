XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A�H��ç��(��n�%�� ���N�!��k�3$�Y,"h�`���zP|��X��M��������Ff�L�u������B7���v�T&?�s/��f��{�� ���QDt,!�uc�;b���	4�2<��Rh.�"�{�:_^��o��fd�<������$�)��zj�'�r���S���gCR~��-��Uo�=�浌�f�q"�̖�j��S��2U.P�7ю]�\!��R4�kbǂc�Y�Ra�ʧ;1J��[A7�:h�?*����:�)DLKO���Xv��"i�����њM!����R~ѽUv1u)����DO���J�#8�2T;��*?e�P\jJ�(�(}�N���B��ww�Z0�#��.;����'u�o;��A�M�!�ˁ���Eg��)F�T)`{�,Z�K����F(^�;N��=��Z\����$�	��/Y��OpaC�g�~偋�Pk�H����3�1 ?�um�\0O�F�L��'�{�B�O��@�/J����+�jH0BBjP�����KK��B��P�@�����+[zy����E��s�ڞR�n-Ⴒ��R��:�� I�f�_`)�k9��0o��.e��2�P��o���×]�}I$�^p�w��2�j�gߛ���(gjآ����
�4[����Tq��/OF+kOBoa.��>��C���q��٘9?�T�f��iǤ���⣶����z���앝t�S-��*���{���P��gXlxVHYEB    fa00    28c0�y��^��F�O1Z�� �&l� !g�Zb!p�r��Jh��g��l�o� �Y\�;2/=�ȟl^�q�Zq��eʽO�j��ĆӍ7���NʏU/w$k�t��3{':���)�D�TÃ�XI�r��PC+e�����j�bJw.�y�.$�g�L��r��O��섚d�ik��ׅ�ڿ��]Ǉe�E��rӐ��|'mK��s"�# J
	WC`9g�&X�j�V����������A_��Y%$���_�^0��Ӓ�G���z^�%���a0�Et�4z���k�}�R���F���!}@)�hƙR$WY�c)Ǌ%,�(
�YTԙb�Jn���8�ߤ�qh������ZYؿr9�9�"-�� 7���EJdNO>�ͭz%���/�>Ԣ<]����������t���O����4 �V��5H
���?Qu[$*7��Ӹ��&�2^���tH*%�H��F��|����-�����hޘ�\ ��n&� %���ѹh��Æ.OIKI�e� Rum~�;/?�̫�Ͱ�O���9��-�Q��ɫ ?#'�"�ƂLJ&�*-G~R2T�}��y����WA�x�cdc���Y��D�B{ߜ�>�5��M*����n�0-����
�5�	�R��"Xtf�����l@��li���R��Q�N�)�� �WgRY�'	h����'`����O�C��r'j �a��Ӻ!�+}T���Lz�+,�'���T���\c��X�fp��+��I�k����o,Ǉ1`�hqFR� w���|����$a.i-��z$�������rf�Fn���i�,�fJe�@|��JRڋ"�d��۸64�&@}1D,}���{�6��<.A$=�V	�#u�Y�\��w��Z�$�$U�@/�O�`ȩ8�uw��l-k���~,\*������$���ؗ�o��a�.���/Ȍa���7]+��{�����絔��FVݽ�b����%��.�@�k[_��(�TV�=����X�����L4q�;g�|rb��\���K=B�ӳLxc�]������@�J����~Fc�=*/( Qii�Ix�n�2�?e��<�&cTɌn���R�����;<���=[[�ko��R��0�MK���~1ه���&���p���?M�4˴���MLn�Oc�
�q'0G_��J/�TXp�˙vU6��X�L�]���3�T�Vt	5C�g�r'i �%B��@Iu[�Y�Ċ�(��o��	��B�r%���1��^p^�D�ʶXaN��6^�v(qQC#|�`����˼u�A�ي'Y����b�rUo�Y��b���F�z�`�$R����_Kgk�����^A/�����-�˺@�N��|4N��"�Y"��F���ى�Y�)]�k�J1��{H�$P�1�%)1�m|ry?C����+B_4���.��0cm��y��Ӭ��Q�:8�>L���	���Da�ˊ��N��]sY/P=��ҪS*�Cn��A��	n���u��n�t{�M��M�`�R��P�~ �������I2�,4H�� �av�м�����+�J(�4�z�Al��
�8��31�j[�X�E���N�G�^܌�#����oCz����*N�w���\�;�J����_i*rě�4X�rBӟ"[jI]���nC�0�2{�g��ɛb0y�S�ި�D���d�$��R������z�{���m4k�5U��k�� ǘf�'2�%b��nD�e?�mv��]q�c��y����X&6Q��=�y"��X)�|�aq�s��/��&~�.A�1q��3�1��SA�rV(�W�Tl{�T��>�WU'�y���>�=6���F����I�E���j��T6�A:�Qĝ�z���?۳6�z���P��oŘ80(w�a��bU�*�Rb}c~O�0��ӷx�}@�C��&�(	�[��	U�EIq��Ag_*	K�4a�zo�W/A�c�է��⚲7�ƅ��s!�a��a��GO^����$�"��; Vm;\bU�k�
B���'�K��l��Fۤ!m��QQ�����B�=�P��5��o������`��ؘ��5:>��ZcWUM�m*~-%F��hj�ʞ��J�ߓ�?�󰝩I�4��O��S,�낶����/*���HcΈ
��VL�ОD��KXD)�r4��3-�@�e
������+��D�,�[�Hôtf�/;�������k��,��x�@���['��;A/�;~#C{g����؝]�7�xɕ���$A���%�>t"���6{�![�6�4j=V�`�I�l�� ܗ'6��m1���%���c��xo�0Q���+��~<��i���Z�_EY]�Bp�fv$X*�s�&_��~2�Q ͫF��|�&�s�ֶuy;V_Pg�乢��O�X��x�eC��LDC�����q�|OA����Y���[���5$�ЏS�!ը�`A+�R�U']'�ѧӇ�ר����&o�S�ɠ��};6��YF&�wT�``�Q���߱�g�~8�nkڧ����K�4�u%�KCQ<����G%����h��Anɧ����o�LҎ�@�Q�^PN�;�pX!�^�
`ZPɰ;˨������ع��`n?5�q�r7<�Z�gB��:c���t�a�*�j��G%��;���B�Ksq��Դ"{f��E.FT9��s�c5�c�]j'`�-v�"L�>�Hi�d�C1|LUϯ4�S�o�I�Ӥ4�ΰ�%���2�8"ɮY�_ӭVG�f���Ǒ S��������_ai{������2O\3�@�|zd��+��ڮ;X�uN��$�L�Z��[Z���d�e�*�x�G�X�1(GEl��/L���)F��AS,��B�]��'��ǫ���/�r;�'���S��	��S9Jx� �7��l��b/���6��,7��ihꭄ�Xd�I���<��@�pWKH���3湽�7�.�8O����Ƞ�R�6����E��T��`�Wp���m��Z80Vq�zi�48# _EWFx�|�FA:Xϼ�Sp�$�u�*�a ���uӻ��h�N����x��F��/
;�������@�^
Q�,��%_��0?��2є�OJ?m��ٟ�'h'��&YGá�z���;��=��C��uU�fKa��k���Z-SV8FT6�0:Ie�C�#eρ1��ҍ��o�XHj��w�̆i��f`��Hj�N���:D4�L?�S��P�Ƃ�� 3	m`��WM��Z�R��}Xs�� �,_��UO]e�ˣx+Gy;/�!]����$X����R	���`�쨥d�k� 9	�L��P~�w5� ���B��71����],N7	�Z1AH�b�F���5o�ɭ�^lkHk����vαe��kJ�������� oE����N3O=2��ʑ��z��",3BYM]W�p�:�n��e�Z>nS�s��%��U5��h&��\�_[���tu���T���ϤKW4����S��C��13�fv�� �� �T8l����b�nZ��o���>�S�[^Z<(�ʒ���}pU#'8�¨u0������.��T��:�c���e)Mw�ԍ����%�g��:K�%���j�/	t4r��y�!M8I"N������(�*��c3�9�9=�zXL��{w�����%���]���ti��X��n��S�pH�Y!i烖>���!����i����+��#vo�(2f�r)�e�4�����/�g��v�SN�"��������L�	��/S�5SZsd(�
�:�̐b�y�/�;טB�JE[E�,[�oZ(��Ml�mM6�V@����gn'mrZ���B����$c�lD9��Gƈ�7EQ�D&�ʘ�'O3ޜ>4T��j-�Ȗw���{�v��sVx�*�#0�����fHpᨌf�5�=��Ձ��\N���>1��#���|�Y4��t0��#]C���C]�̟AH&a�jRQ��UO
��Mv�4{���0�
��[�ȐȂBvtw�q��� �r�tE&��^ID�o�R�4Yr�P��i��o�y�2�'����z�\���W,��m}W	 �_g����i��^h����]R5L��U|%%�f�d7d1�,�DL=��{Z�';<��ANp��>	���`���rq4UNsiX1UBKYhSfHz�`o�/���*��m���"D�ً�6b��g�qK4�� �2i��� z����Ο�|��2�~k��*W܃�n�-��%�A��ڈdHA0�ʦ�r��an;{U����K�oN��4<j�)����ۣ� b_�3�@(�'hC*l*��Q�Ҙ���^�]��Y��(Q�~�H���i�4E��3��ȏ�^��y>��d�+�٠[�ꢃV�x�iA����a�:b�95� �)�'��CDߵ���Vrο{���Oy1d/���u��p��$�F�ξC��p��t!����`w����!�!��j�3�$Sx]�)��;��*5:_��[���WAt�ɝg�@�-���c$�J��kN}cE���"w����I���%��3Ĉ!�F���� �G�u@�d��.ě�,7D�ch�,%��:@�}(��8"rm�{�a�m� L8B�Z�=#0�V��������Y*��M�D�d��3T�#
�h^�G�����8���k4Q�^ܥ{���OG~�K����>0u���\�y:L �vS<Ć���Φ�8�T�dr�	<[�H��&ш�uNHoi���)��sܐ��7���������h�dA�l-������s4�{���"nwL�Rv���P�ȱY,�3�w/����X���R����a@� �q|����~�)Iߠ7 ���e��8קA���*XXC�b���GΌ��O�&���O�/�0t�����O��ڢ���}�;��b`��B�/���d�<_�kνg3#]��}sލV�Ҫ\
�{b̟�S�x�ML��A�ؚ/}��N�L,Zb��ם,�1�3�I*'���SA�i5�`G�*��� ���b�_I��{�C\�.���R�c�%�e����ib#�&8����?�W�2��ژ��0>�&����0���u���Q}9}BAn��R�J�s>��If���f�(��-����t����Պ�XN���fOf�S��]w�����
�GE��#ՙf�c��b��٩T��=�̥ ��N�����LLw\i֤}>}���;7��x��n�{��N�z�lg煨D*�ȪK���9�(0�\���m���#�W�c,zh9S�
�6�H�̈́MEF��]�k B�I�1?"H$���6Sm�� ���$3Y8���R�nc��R�eZ�ĜV��=��p�L���\�Mpi���u�HO�X��gΟA#���˛���׽�8^E_؛"n�f�����Lf8{���V���@��<̋˖]�������i��Ǯ���+�~�����|8��tmS��w�	u�6>0���Ax-�y>Mi@�%�?I$w�@Ǻi�?�*kq���#��Gm����(�K}q2�j��g�����:�^ }H%7B�"�(#]v\�I�1VY�Dj �¤	��>��X�,�m�$]U��cs�C��D�\�yFQ���̟,A?�*�%�F7�Q��2�����5r{�S���	�� 1zկE��Q0!�ZW��G�3RM��H<VӰ�s�mf�x�!�;�آLzh�A#l�����t��
p�������l���t1Ƴ}(#h����m&j�<v�,ʹ�/���;�C9��p�[*?�\�F�p�iO��_vY�TB��%ᜡ�<����u��q+㳰^�.�0��y7��w�#�C`���?�*|<mw)�u8T�URf{Ϛ�\�/�i��k>G����>jJlXM�<*Q6b�*�5��i[��R��ϝ�;��	v���r	UXS鬠��3�y϶71n�/����>��'�<��KS�_�E;<�xY��t�F�I�z?"�^[-F��_��/J�� �^9�d�H���g����C���A�g$���}P�Jm��1a�h|�#���Y�я��,n6av�K�
Є�+yhj�+�t�� �;�� �oS�^X�l��{`�Q#đe���4�!�>�`��D���
z1D�4���H�132�,���S����s���Xht�%6���~/Z�]b���t����L\�� 6O�BM��m쇰E?�Azį�v�zF��O��c\$�@9�,0��p��D&�)]\��><�ӂ��������b�ޯt��X�gb�lJ�J��)�L�K��A�A��c8�A"d ���6���J�� G�[q2&�̬���ݙ��*pܲ��Z� /�!��ڢ/ï��9D#�'|�;s�`�F��D���\�����y\2��r���m�|�!�&��v֬�4��7N�D��ٔ䶀Z���fD;lRS��Ʋ\2���K�9�Y�B@��g>T���=*�u�3z���Ӛ�Ai��+Qj�#��͕�z}E�"����7N#��z'E�tzq;)|�f4��"ߩe�_Q1� �*;s��>���	�W˚B��(1��s�V�kWir��`��9N91���i=�� � �H�ۯ�}�e$����Ow��Kk5l�ô5��?������-H�"e�o��D���`��R�^�����h�/0�H<�'Y��|�k�a���Ĥ	�C���aK%��D���x��o�Y^�n{�ʼ�%[W�<p���S� ~!$6%(��ʪpk��5�h5�#h<#%������#M���H��>�5���o����d�G������s�P�MR���'I��v9_�;�t*VU@�8#*�֕��p��L���$Ŵ�5���u��k�.z�(�^a hCX�g��d��m9u$�9��F����rz)�/��[���ӑa����b�?(�C�:��wj�HhH�0?"NG�'07��~�x�N�
�q�
�(�Ѝ$?
;ЉD�Q�y��Kj)��gM�����0�QS<H�1�)�SB��G�U�3�S!����f Ї|���20Ј�������Gh��Co���'�i�jxm�.!�:Y[�;V����M�ƣ��s��7@��K�cu�R|$x=D"b����4�$�s�m�HT��.���מ�F��>bo�'���vT�����<}DW���6b�>|Α���%M$�dD��n�~�;�,I���rɦ�IǦ�Ѝ�oI��ϗ�����Ѫ�H5����C�i^L�r�Rc�?u�.W�zJ]?[R��O��_2?��5�*eU���l"����A�k��dL�.[��D�X������P�t����l��U�������	J7K�U)e�Ѽn��� +Q��"-���HK#{=�)�,� ����f���{X�v`�S�5V�մ��9;]Z�+�3�t���Gn��٢��~n�Y��$�/S��]JO���͗*.�|�j8�ΰ a�k��4,V��qv����*�[���ĉ;>@w��D�B���ҳ�Z^r���^���H�^���xs�	�οk}�UIm�K���ч������g��Ţ�G�i����.����y���Q����a����)�b�[�%����[w��F��W>���ʕfx�S���fN���7�FB��[��*?�.s�s|�� g��]�'������A���@�K�=�G�1ߨ}���Os�ss�,����`$C)D��M����¥|k�2��2u�����3ѣ���w�����,�f�I-ȕߓM03�cm����������N%�� :�;�~ s��r�N��~k.ۃ"��1����e �b��1@���?צ�4��i&����%E�Ã��S=jO^,s��};��jD[g^�s�J����uX�G]�Y��~�6��od�L}�Φ8�J� �qp�C�*Y�}���>#U�㼑{Z�dO;�l�p��i	$Ie��s3��H�k_0DI4�&sSZ�}�ʪ���+�˒0�Gpv=[��1��q�2��F{�Rx"��^����>F-+&:N:�~�d�M%Y��FC�B�ډ�]��м!���]�D9"�d+r�b�I�ng�O�r�NZ�D�m���}���� ����d%��C`��u�+��HH���\���kW`fĎ��k8��H�K $������F�(���lv�����{:�,���L�TL�(z�!��3j�E:�C9���Xu��@'��$���-���'��/�ٓ
�|(P�|'��������zf O%��Ԣ���H2Iߪ�_:;"�upk����Nz�(o`TN}T�vc6�#���P��2�9�.?�Id�1���{�T�4�[�b�j�X�|vIO:����+��'4{�������#x�$#�����,�oaZ�x\O%u�e{��B�����㮛u�i��ͤ�OF�.���#1�8���|�
[ݮ�l������'�S�2>.W�R�z��m���W�0��	is�ظxFK$�Y[�ܦ&�#~�I|� e�`
�9��{��0S`�!��x��%��
?���W��ayE!*3�(�OY�A�؆�̂�+_���eo�N��_�4�.^^ ڜ����ah� {�T��Z٭f��5���D8p���Ca��w�!��-�I��sP��e���I�wx���D��v=�5δ�s�9�S֒���m�.l�f'LRrl�Q��ty���A�K
�7�.E$�ni�H[�'��NE�w�AC��jD|u've:Z\��<~d���t�"Rd~��3Pu�#��Oז޸�p[��pZl����7nU?+�<@��_�����@�&�Ç���L�{'�O�7��S�	Ud(�4��#�HБ��^��a^�.Ԭ�:o��n�����t�8V��^�7����dR�1>�����hzs%��{#��[}T_�>D�BT���X4&;��,r�J�vQ6��{�K�?ʗ�P�Y�ah��}A6?�j���g�Dq5
�E��u��h����4��|��}s�՘O:d�L�Q�o���I�������Ԋ��1*�k#)1��-��2ʋ�$��0������5���#��[{_f���w#E=��\&�±j���~�(ΧC������Q��b����Ұ�58��O�{�����ė/����X���D2�w�{���"����׌�R���V�
����l�>2e�Z���F2HC��$C���며�N�P��̙6;�Y_�u~�eI��N��h�X�V��*o{Ga�[놝qEh�(�4V��C��y�> A`�o�6ð� ��{�Dp�SY�#����Zf��ۚH+���d�~�O��F��x,�i�Ĕl,��t�s�\��v|��4Ҳ�I���sS��n����h�"E��������ܰ��&�:
%`,���n&^ B��bqn%}�'KPޡ����UC��΀�W�p�dgQ�Nȫ�L���UT8�m�w���Wsa���X�$Ho2�?�������	0�B�	���T���E�lp�aR��/�_lfyE��{ ��!��ߐ�*�����K�I*�� DN��,3٤}����q�@��e��)s��?�н�컮��߅�6����Yw��M���iLتK�*B��#��%�Re�F�޺�I̹��/ؙYgjˋ*��c�{3�LN���cN�H%�6�.@G���ו5��ϙ��x833����\!���^���_A�ix�N����;m,/ ��x�qSk$AU�
͌��U`R��ݚޙ	�ז�^��tƗ<d��[��1�k�\�i
�9��b6ܗc�&Ț�#wRC�$D��x3\��숹�qY,[]n�>��4���6��� Y�4��E�ֳ������g��NH�)�bmƷ���R���@��?ܮ!��Wi��h�8�5�J��j(S4�i�!�M	���P}_�0�Ab��!��f?����m�xkw-�X��J�6�,�a���9���K��%֙M���!�
�ې��"k�*>�ntg���ҽ�xp��I��rq����kn�i8�#�ߢ�D��A����/2��z+�I�(�`�Ԥr�� �Pz�}$I�MH������ݮZ�:�y�G�:&8�9᫢B��k�t!�HzG�I-Zkt%M��Y|yֈ�"�惍�m���%	���y���7[@�(����^�)�r��2�v�M�;WNӬp��o�R&_Uڙ����34J�k�E�Jp��e
�!�+$�aBTNSE^J�*[�HXlxVHYEB     896     280��+4�J��n(&��j�kt�Gǈ��Z;2̵ ��&*�4>�9�69`�
�8�K�n��=w2,9D�/2�6�
�Q�1kA��P�ƙ�b���ﾷ#W���Eq�R>6���_�jM���#	�h ����N��"�f���N�Qo�P-Qfѹ5�A?�YZ>_�}t>
���,�3"�
:�l@bW�u�P���	�v�>�	m�H�9�M���h0��AC��)^	w�>��6����Ҩ�/�\a2���^�R������?���Ҝ�)X?��G�7�f��](���\B�	�ͦC\,5�kJ���I�._�:��Z�.��{^�>S]?Ps����h��z��Y�r���5lQV�����5r�R-Q�x��b�@������ɠ �/Z_PW$׊���&y���~c9��!�	�ф���Y�iX���#\�`Y��s�ը������2���; ���6FE�v:z�3熤@m�o�ԃ�Ga.������N�׭���\�6��q0vE���ᝠ��45�ZY�<y���ŷ����'��]�w��� ��ExoKY�%�4�Z����avm��λ�7�5�Pcm]t�l�1hX�-��.��5�M@��2��R��M