XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��c�)b��+_���Q��.��}�_޹������m����Ң�,z�Hp{8���lIkq�����.�+j�Ĳ^#h�y%�I�y��H�r|�Qіa�x�݌���?:d���g�dڒ��b-O׫\�sK���SD=�5]~����u;k
�|K��K���\�\�hc�#f�b��n43Ӄ0 #�}�@�s��۱�a�����O����� #�Qv�3@��������{���Մ+ �sB�7�k�Y$|���H� �nP%�H����S��v� u~�8�EZ����Ӭ�I9H+�λI�����+7���m*Iau0R��|�^�N+�.����S:����Y�b�4+'Xkm*_�r�:�9!�}�{��#��#�v��}�G���hȅ`�[k�����<�n�{�CX�ρ%�H�����ԑ��3a�N�"�&j��Y�C:���u6b�P���dlz�dSp��3[�G����2M���NM]X�-�)�[����r�����;:?.�{���8-J1�y�v#�E����~<JDT��K�� �Ն�ht�2VA�p�Y2��y���@������/�j])��^A�� �����d�n��9�M��j��;O���ٶ���S��=���/i�{����%R� O��ӱs;zBh����TBJUy�����
~��Q8�!�*[[�q��z_%`n	����C�[#�o1ȥ3
�OM	$a�zlD� �N��Lk�&���G�Ig>�he�(5XlxVHYEB    c763    2600l�X���5 ��:-x ��[$��TdId>�)�+�:`Y˞�2š��I��_�d����
f�z��p���L����J�"�Vk�
�إ�67�lK�X��Uk��ùގl��0/賁kd�����xM�N��]���eh�[�%
Y���|��Gh�+�/�W%0��M�$2���:LTTM�-��j�1jac��3��ٳd��SZ}�q�4�l�	��ʵA�9˲��Ԫt�K>s+,����陼���ި�W�w��D�g�iX��ӃA�z�@b��Ɣ����L[[�Q�*��C	�j
���h����*c���`�泤�3�ý:��G�\�a�'�R��ܨ���zZ�݅��n	*��_�)D$�JQ��O���K �9�d�0��L�gp�g���2�6���57�a���"����H9�6G�z:;�4Z߮��Y6@M��׏>P�;�$�����G��� �;D�kF�-���h���KT/�#W����gn��C9���
~Ĕ�ڽ�B#���r͘*�6�\z�k?F�P�6�?��fw(�f �%D�>��(�WW��̡�6C�H�0M��BO����q�i�X�����_8�l7�!=����m���*�4��h�`
`A􄳭^P���*?��(��;�9�Ö́-&&��p-�MUѴ�u�4�bBY]y	,Ԁ�Z�d���rUyx!�d�¾|�"߄���\e���S=��HЅf��.z 8��B�C�fDN��Ȥ��J�l`��Aߓ��7[��֩	?9�>���woD�n�	٤t�7(z���ȩ���ORu�+���}9ݽ��j��9��x��a��H�V�yd�Y㓒�h������Na"H�S&э�'�<��7,�(�T�C�+�d4��X�����	Yj���2q�2g������ݔ�,I�,cX ��~4���bߕ]� �2QY�dV�<_u�V5��AD�a=?E!(��6�yj`৯Ink�}<~p�_>s/>^���d�{�y�T^ԅ�Av�C{)q]	:�
�-��ܹ��Qo楟-����*K?���h'rЅ���%LIiQ�2���߈�۞i䲯*�9Dt��J��O�v:�.��Kd!�vA�]1�8hʎH���#K�NSK�%��xb�ի��M��� ��Zf���'�Y��ehp�����yv�������?g��5��D� '�v��\:���sh3�2[�N�"�a�w�����F�<TF��ѭH ���7V �ڊ��IBȇg,��F9ݺ҂�΢S]J-R��E� r�6�2�!.�g���2����C��U�����c=c5t���U�g�-�� t������ب]-8��K8H��Zb���V�1o�^���h�����㔩[l�E�}-9�,n�*|ȴ�k�Tc9�N����� ��J̧� Ӕ��)=8R�W	�xBi�����d��/�\�S��q��F�ʐ����K+@��R�Vՙ}���G|0ɔ�p�Ux��д��XV��.��Ti��gwI�sK��W�1խ�@���繓�ƽ�[�B��]
�D�{��>o4Q17ۦ�H<Fx����X
�T9�:��0#���s3y.�+����5��9�n�B^�&Eg̉��*��;��r��b2׊9C�/��U=��M#~��,��P���T.�_H�T�7�Җ�x�7D�o:��r�nYY:�Ў�D�\��tx�D\�_��5�9����LOZ�/��|^5��>���SC&8rzg��&��e~����=�_� �t��hj/����W�8lFvh9�OB��Ǽ��S�Z(�TIhVԶ�#(�{�l��	��r&�����²���Q�~���#�V��Q�)��4�����S���l�y'~K�<ٵirG�7�ig���'lfU$��g	���v���齸�B�
EȘ�4*�-��)�`,�^����[K���@ ��+%��1\�m��S̜FvN��bܐ��i��Ωy�?�����e���zg5[o��ձR�����T��4{G�kT����k���U��l�9Q�}�����x�ia.�-s`�H 4b��e:��}G^��y�3�U�cD�Z��l��\�ݔa*�������<�yiL)p�/�����~��I�{A}knX��t� �k}�ڨ"û>�'`�k���i~Y���$��*��_U�	y~E}0=L�O����F.!�>���k��P��@�"=�8������s��,��N$�)
O�f�Q��~���!J'g��$�m�0rL������y��>����K�V�B�W�ψ ]�kz��3����4�P�{'H��@�I��Йt���J���� M��_p�G�^\��@��e�L�_;B�Sga��\��|'�/k�.����d.~�u5�4u9W���V�S<����,Q}NI��t��m��X�X�z�ڲ�����Bƌ'>Q�xf�"�4�#]	�6K��6�`dA<*]K�[��k�q}��X���ܲݾ��ڿ�3.�	5c�Hν��5�����`]�+1}�QJ@+f�H��"
�<l���?�<�Ց�O<6ω��7WJWp�Ң��A¥���2K]��M>�T��
̃�@�������>���!eg��uF���B/v�����h�Q��4[�k�BI��[ӶqZ$z��Y0jE�� ��W�NU5̪y�;���FAڄ�&�o��ۿ�"��q�K�*�E�ў�_ ���7ƅ�Iz��c ��p~��.c�j[��?l�)��z�.[�4h�}Y/b�ٕ������R�W��v�#����	����/������=a��5}�U>�"�/���B�|��,
�)Xk1������x�6c[t\x'��\����Ԓ!F����gE±������rg����zи/�F�l�XDl�}n*֌�5�ϝ�X���X.6����gF�av�ϝ5��ŶϺ���X>�B�.���Ԓi��]��B�G�=��GXm +���PL�tv���%n�\|�Ǟ��u*��×��_j��ҙ}1��<߯���/�}��9�p��\�i~"|���?o���W�T��U"e\��=XiO���
sK���b��Ť$�&��@��`J:��A�`�-^��B,}vE�T��}�8��:p#���!���E5d��M�3ສ,��t����m�P�%����2�Fx�m1��{pDnj���u�^K�д�M�V~��˒'�FD>Ӄݸɬ��;�,��:��8֯mR�����aU-r�^^��3�.�ދ|���O~�r)�yJ�`{�jc G��a�d��Q��%�����h'����4~Fb����5M�{�}����!���퀨ވm�*�Zʴ��pnnN�3]�<��5@�ʭ'WyU�}��BZ�y�N�P�؏mN}mvf��:G,��4��L�^5oB��|�r��`o@�����*�&�%|H��PY����zd�Jc�E��1m�6�l��y�1�Q��4�R�ܑ�₳c�����n>�E1� 2pg���2�1_L���Rpj�0�U�����=�Fɢ�W��T�f�52�.�q5C���Gd�iv!_�v��\u�h���@�㆓ �H��7���θq�ۊA�2������%AYЕ�BW��yW'my�i�qp`ɜ�g}�'(P��n[n��>��>Tb�p�bCj�ѻ�<+$P�O�7;����p&�;��Ӕ�1��E	�v�W�;��9� p�3鵜{�������jM��#d�D
ʙ��R�G�Vm��eE���W�u���侗�����d	y�&zw�a��^�n�"Ja\￭����\�;��4蹶���cܩ�.wY/�٪؉�&z��F���52�����f����I���*���mS��-a�]Q���+��J� ��{�5���;��a����!��s���ͲT';��2���;-ik�@����	��(q��� ٴ�B�-^0}��u�\�S��^hh���I-��VA�0g#��jF�Q�$��|,1���3V�l��-RN��TB�`?D���RI����������,�]O����j�����{d��q�L.�c����w|+��ɂ����,X(ɴ}�W�<� �a�q'	��J��pG������:�6r���^��"%F��gAxA"�-ł�?4P�T��>?W�W#�g�kY�b4<Gh]86�`D��i�Z(���E  P=H>��0&%�2��Bv��d�� ��?T���6��h�AaK���[�Z�;�d�P�=%S�	U�C�<�w�Hk�ж_L�lB�h����jp�-|�bqRK�~��g/0"�(���`2r�~8P���L�'1@�����%m��~�_��7��L
�?���	����㍦Hx��@�����p��챝��]72���}	��K8	�0�^Q�f�a��H��a'��E^߀Y��c�G'q>��4Sf���L8����!�!ƛ�@����3Z7�t�������p���L#� ����NJ+�����3{�t�ʥ��.{j�ݝ��3���Om�P����w����5˺;�3�0����c�XBG�Q�J֟�lm��vQ�9Hn�0��w�5 %�F�ذ�x�B��/tJ�����x�lx�L�0��q\2���P�A:^G�j�h1�3F��X
�L��+���py����+�w�(��F*�Zx�2�O;�!	\ل3N��,��j���Q[1�,*|�]Y�k�O�+�|1��]��B�v���i��o�yUV┅�oN,%�6�I�v����Sd��e5�t�Ќ
W��B��؀�::�����%;��msӟU�+$�Q����2���hC��ۡ�[(둪$��t�j��hr�c-�,������ß�=$�!<M����	|[�_N�o,�,����[e�}Ա/$*$��|���`���e�Ò��(-��#����຀�̓��SU!�*̜� 	(�M�Iג{�K��fz�f��7�Ԁ�8KTV{����*u��N��4�"��T��'$^�pZ|��5z@��~V�)���*GJC��	8���1K?E���8K;���'oJ�zQz���YuvcQ:��x߬�aRv��YS7�� W&���@<"��G.�/�;|#�x�D�K2��J�{�EN{D�ĝ�c�T��Z�Wh�����ih�Qkd�Q�5�2w�D�I� �Ŋ;΃z����"�������ec�e_篋13�]ې�����,��L��O˧�<ivU��Ԏ��}l����z���/5U�i�o,e�E�Z�s�t����U����L3I7;噀�L)\�p� Ž���9j�g9y��f���w��)���$��R��t���n ���l =dnL�S��i����"W]}�/�XI�3v�,�X4<��)nK'@���y$PG;%�Cv��8�fSV{ќ������[�BhIF]����6�A5aZ�1̫�V`������\�cp�Ҭi�������Q2N�gA���]��I'l����H������p�:�7:cb�]ѥ.7Y��?~ե�w��p��R>ƛ�W�b�c�Ē��W���rn����n�L�0��-���a��=�]��H����X�M�*VØ��1,�1c�l/s���K��d�˸�1��$����X��]��չ�k�BP F�fՁ,�$��_Ѧڐ&.�0{�ܸ?~�������6#�!-u�\��t�)խE�}p.�I� j-��@YT��VF*��JN���Pr����{����e�8�ѨTt~�+�ĜH���{��9�n�R��>���#���1�x�D��P����$�ڸ *�����ZZ�39ᔞ-*�s���<�$�&b&-\�G�o�;�%83iZ~Bg�_7�Odrá�>���n.�+b/k�%�V������x�=4z2� �w�����Hj�#���n�&)�˸��A�'�<�$vd�i��oճ����u�
�o�Est� O�g0XD=6E[6U�׎Hi0�A���7�H���B���Dd��A��C@�Ze�_�̄��u�iҹ����A��W��0u%�{�WEEs3ɮLoJ��ys��D8V�F�gXn�ؾ���Gٯ*�G��pcH�5��8F�}�<�,-�e���*�F/�q�A�9
$��&����K]�`�]_��SWv�t�sx������oF��
�������=2$������S+�#�9��U��{�g�57y+��ARU��wRq����*�e�y��셽��Qͻ\�\����y��=��_��:u48��I4B�n���t0����c�>*tmd/�s��
[�d@��qy���~w�X}Ƶ��Cw��7�_*�G&�yB�u����I U�K�8qOFir)b�c���u�����;�k�s��s*B�u3)żhY��|ji�rP��ƮpneƤ5����l\�����S&��<Q���W��%Y����.�E�Ѫ7���p�2�HX��4|]ԃ���D�~繸Ĉ�-1^���16�;"�Nf����:-{q�P��Ɋ)/�e<I՗����ƁUޓ�,��m���ۛy��$�<)��R��������X��������w����`��=b���;�~���$@e�b|#�.e*$�[S��VR*�OnSܴٸ�x�m��Ql�Ma���,��;5�q�*��=!�I�p[��~�����z;�p�il���
�O+bv��JSl��;~d��H+?}i�I��󝃦O�X5�G�a�'UMw�� 	���AR	�dy+v�>]��b����EJ�R!oƟ�D�r��ِˁ��'O�њ
M�V���l �H�1�����6��.�j`d�e�K#�O����ש���`� ���4XU������fU㪊ɀķ��9&.�N���\c��3f89�kMb}��m�#,��Q3�n�æX���hno@��A�j�t���:��d�˶�e���a��_j�w�N��c�*;���u\���	��w��=��>���� Ź�p��)�a'��X1����,�d��o�#�!�-K���>#�+:X�M5�~W��j1��!��Y���_	��q�G�|»�Ȓ�p�Ԋ����}����}�\�����YoV�����Gz�\j�/Ɠ��F%t jN��&݉�y\��Z4&�oU�v��>}�{���=��/&��)|�z����zw��(�������ӠpC`u�>�)�����G�����ӀE�<��;���5[�F�ԉ6�,����W��h�Z���6?��هHc���z�+vq��k���6�xosN���"�����I�J�;q5�*u�c`�%9n;{�@Ҹ8��ﭜ!R�ԂSZ�㑓�0��<�ӊ$�^��v!�X�����e|t�/-Z��e�̬|$�wm�""=;&D������m[�AC��,�5����CA��74h�1���|�*u0&tÕ)��|[�KU8�1����X�Z'��3�L�#tF���b1�8�ڔ���LjD�j�ShA��ÜIIy�K&����{���3��^������8�p� $]e�Qg�F>�J�MU�S.���m�H�+�8oB�/�j$��p|�8x�JL��L�ݾ�x�e#f��s�j���2{�)���U�g��bV�W���3��|��T��K�	@��$X�į����;���nJ�v{�H���wEd��e�4cl�\z^�J�,sS������C��Ta��)��wk�>ži�!��t�ݭ����:�0.YgL�F�T�w�j-���\9 �6�ѐ�~�M�2���#�a},���#��!3���72f�����H{� ��C�_�����28��}(��T�(�#~�pS��tá\��C�x�zaEcj����b��q���c��wA	7�
d#9�}�;@�z.�r����!�i����Ъ�^��L���@
�n��# �6��}	���)(��������p��r��M�<���9AF�ӇĕiB[�p���M�A�ՃԄ-�p��d���ı�Ѭ1��<o���Zt�r��t`i��_)b���(�w������N
�e�l	�2/��q|a$��[S'��q��'��;�	QYߋr�7�5�\� �7���'}Y�
���W���T�ڳ�JIj�kio���Q?�X�Q���f(�nEA��jH^�DP�I6��A�wQ�DD����a�c�m�;�!��qf�ݺ��,Q<EKF_�? ⁥u�F�4���x�G酹����	.�9o���(�8��#�4�Ok�rb��	�b���P���c�.z����� Z��1"�,[~�f_#&b����W4<܃�Ճ*k����4@i[��7S��9z�%����:B"���*>b�R��䃰�ي��Vr�ݪ�?Og:� 7ԫ�M�T����EE�fMKw��b2�c���L�vh;�յ�C�"�mߦ�"y�����[�wSq?i���QH&��3�� ,��EyJ܎���o��J�OhRYfThr��v�/��\�ym搔<k��qh+���@xvs��`TI�!� ��T�ކ݊�]���T1q ������,=��c0�	�-l�v�χ����������P����먍{��3n�# �Y��8L�X��"e*ڠ�,�5
6Ɩsv�1�[6�!�Z�q�Ӿ�X���9t�C��ۋ�*}����U�`���:��,����)������c�bՈ������K�g���l�� k�9/�'���,����$ٶ즈�$}�!r�s��j��#�_�'���'c�o�Ҡ� 5Z��i�9�'7=�!��/}��ȫ����������;�C�t�0�~�c�Id���x��jim�z!���^����	Vpmа��ۅ�I�	���=eNI�����ɂʼj�R�`:�Ś��)*nQ��� ��\|ٕ�"���,�� MĒr���"ɧ'��{��g��w54>�� Bq�6�8v�9�
Egﺍ42Y�a�H�sB`�u��v�<I��~���+M�2BB�����#����_����N��'�=��xH?^�{Ӝ fs��cX���2>	ס�	͘u���M��jD7�'�Ç��L^꒧����ɋ7-��rZl���ӑ�DH�W8hE��*�oY]u���&t�4����M�Bf��^d�uV���[X,���o��ތG��b�[?�8�ގ��T�4K\����t59��FAK.q����4�#�ė�ޤR�^5#omC��=��:C�,a	���r
j`ܕ�PGYi�Ã��dx.Q�]��p�������t�A�6$��%`n�����\E�� W�œ-��lT�e5�3��(�>��WE�B3�oA�Q|8^k�����1}��)_�����w�Q�P�W�
�]{�,m���۵��K�DEC���,�<v94X>�1j�-BXo��}f�eU����<��/�bid��������tr9w4�1������d֤����*��9[b�RX�UY /�O8�nfU� ��I���h\�"�ڶP��/��9��_��<V�k���'�bԻORKڏ��������lZ���Pz�Z2"�A��qm]١+D?='}d�ͥ}���