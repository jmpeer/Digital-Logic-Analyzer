XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��H��Q]tNUj�1�"2EL�W���Z�qug�lc�:.�5�yp�F�r�?��r�/pPt�2[3�a�ģ*�H�0���~:Q[&~#�:��*q��V`A��݄R�4���3>�Pr�F���w�� ̓�?���p:��2����j7m����)�����Dw���b��2��Nf�<3e4��Q��o��$��S� �S�C�hպ�ǟC�0�}��K�\\�Ҥ�e�û&����7�2A�J��q�?���W$��#:�5�<0[o�16�}T.�[b0m1�R�u��T�Ad������Y`�^��]�;bT}0K�PZ��|���Geq��T~�Q/X�~jA:3���{E�~��Oe�^�]+h&�@_���8_�Q�&X����.3�^���1>h��(e��k)-�x������0�Zdb� �@Q�@0{w�ēl���~�j�=�D��2��˺5.�������K�M~�v:I�N��/�=1�x��*�g\���t��m��i����J��l'��P��^m������4���ô!�c�ܸ:���{�%��� ��	A�<����j���g��<Gl9Xw�}���ť�8@�JR�z�/���������o?i���"�1���_���)8Ǧ�L�{�ḱ��SIj�����Z�8�w%��/�,~����bq��!��Ji��ڸ�7��웏7
W��OO��I���U9~�ZD�Q��!6����I��NHU2W[��KńJ-�Ы �sj_��&XlxVHYEB    33bd     c90�cS���N@�e��v\���k��6+sτRU�3�s>�w��쏐/v
2��ڗ��!H3^niL���s��9���0M_:4}��4�3��|���fd����-kQ���ĚH�A��Ī��*�%�?O�A����ˡz�� 0Iw�M�c��E����ǿ�/���1�B�	�\'9P*
�E�4�|O^�yds������J�.R��bՋHa���4��DJ��GU�MBf�U�~�����>#\�[��	��P����'^o<Q�g�cM�$&�􆄴>ѿ��C�_�b[��Zd��WFT- �$T�铤H�˛�X�W�)�-="�u�/��#WK1��N������K�L'"���s�zz��|�&��P�St��M�Bm�զ�vs���	Z<.�Xm�-Rttq�������Z�-g<6�� �7���$�~f��mՐ��:{t��@�-���T`6JJیH�߽w;�io���g7���N�ǅ��Bq�Fd��}A�("�K���!�i�ΓԊ没?���8r�m��gվ&y�V���h�p��io���hHM��&�懠���CY�ִQ$ �ԃ��z�0�%��Q�?��Q�4�Y�|J�����`����]n���_R,�ξs���[�@�Z[`��g�9��]/s�Q��u��
A�N0(��'�֜ރ �v�7�U���a�-w$" 2h�s�Hm��i����n�/~#�:l��]��W���9}u5�ٚ%�_q��O��{G�a�B���B����@IA����\(��%k����IŠ��fT���j�����l��w1ok�-��7A!2�����MC��J��uz�Z�~Q]!Z)X1t��k���T�	.��+J�I�g�M�*�+jI��zΕ�!\q�8ӆ�#�����N�S��b��V��+HQAI�ùF���۹�M�j��m&{��ɴ�Q���w˝�3Y��t��{�}Dl��c��f���v[��l����/��V���iW4H_j�h;Lc���o!F���п5���	w+:�)}��Q�7�[���]�����(��[Qg�5�#�� 0ϴ�E�������WT��l������]�W��j���ǎdЂ�oz�7p�DP��P��#4��?M� $�T��\u�!�Y���s؄����o��В\�:x�]�P�tG�֚B��P��a�ƅ��A�I���lA�BֈhG�Mf���k�g�_��0L�(a��b�q� ;qd�̾TT��y�(A�Ќ��V���t��5�0��ٶB�DOgj�8�̼�����_��:]�Q����Q-���)6+X�_�?D�3�%��VL�
AUo� k�)l�Dv�ry� ��)���Z7��p����>�F��,��95�su6���s;$f���Q�۩��د�N��b.�c���Ffi��|�I��B��:q����j[�W2@�Z`<ѐ��;#HvYp����{T�]�s�5�J�h/��,�2.��{mf�C�T=�o�+�Cҁ��;g��$}�	ro�n�А7igq1.���St�,AfS��[a;�E��D��@e���_2 ��Գty�`�$s�
B�Ξ*���i`
^Ϥ#��{�lխ��@k�l صX��q�-��9�h��W$5E�I�~�b�%�y|��%�K2��c�*[�B���aim>	���oN
���{6�e�5N�R��I��k�"!��Pu{݈C,��(��;F��=�����ӄ�"���A�!F�[���z��-��V��..��_�/�w�쟊�N��K�������&��؜o��=6�p�C�f��� 7��
@J{Қ��u骺��p��M�o|�3�����}w̡v< �D��k�[@HB�L�KT:9���=� ���9`�օ��9��}'�L)~~c���r�J�ĝ�~���텱�Y*�["���6��C���A���o����Ke�h��"���,��&fTo�a�4R~T�k���s��f� �U�}=���� �?U%���!A摶�ki��t���.��=x	���O�a��$���MjN�� {���Ϸ]^xGX��=��������RE�0V�]۠W�3P��=R����Mmi�r�I���1���!�R߷c߽φ�ID(�S	l�0W=ezDsG�giA5f��0̤�����pqe	s��$�[������v�1� f��h��w��@��b��{���������Ϣ�褚��(��Nä~���"ar����r���׹KBh��@nQ{BdgQ����d����� �]'(��q9pfVY�lN�)�k��tr[Ѵ,}��F���i��þ�CcM�0m���w��BĆ���u_�3}�����f���	��.Ew�UJ�K��]ܐ���%P1�dK;����R.����a���B<�cr�	�FJ_v��X���O�#d@�vC-��$
遢��G2�$��Ϛ�WY#��`egp.E�CD�q��b�Z����I��eX�+5C<9m�Y�=�41�bKˀ���˹�;rHE*��5(�6�H|A�߫J �`�R�sv4�`?K��0������Kˁ6�]��<����zKR�b�Z#+�����^A���O�;�[(6�/C�����O_����}Ԭ=�����7Y[Щ)�%X�(�?����tJB���b� j��L��.*P� P�-���G�� pr	�	��l�@.�&��|�F��͆������\���]!Y�wj���{�}S�ӗ��U�Z��qV�����B��P=ߵfb�G��$AUK*X�%�7���Pd���M�ܾdL]��!3�Ѳ@�����@MfS�´�:�<�����T���[�ڑ�?��X�:����P��Q����F#�=y���]�Ђ��)�-�Y&�wi��m��{���<q��+'u��+�/&<�e��Վ%]�}=t�^rQB��N٩q���C��_F�\;V̞Fd�
N���/�EHowr�+K���l��_�2���}n����)ה��K���ن2K*<�k����>�k����q�>�h��3�1h(��~s�w��$��z=Usc��ٶI�S;��,Č^"��	U��u��a|%0 w�vPs(�Ж��������c�7It{xf{୓௝A�y��3���b�홫��|bX