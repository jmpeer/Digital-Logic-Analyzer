XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��j��ʇo��Â]�*w���f�E4���+��݁O���u����u���~��`�״��rz~͓�ա`cRd2:��-C�.S�U��S�
�@F[Y����-U�����֯�|T*C�z��>����;6A�pl%�����K��/��Jɀ&�_ ���ʘ�O��^;`1�P�08P���׳ȴ�0�SO�Yv��4�K��-�4�e�'@�����{Z`�Y^
�Ywqx�0��9��*�3Z�f�Y�{�	sя�&�@U�O�!�k�ݙ��D.��6/�ˊ�[�)�s��9ej���h}����x]rر��
����m����la��pφ�!�	��&����۰�������L��
�{�&�u��κ�H��#���u��+���cXq4"L�� ��^$#�]��2Vx۰�;i't��v)��p�8�_��w���oN���S]o�?�~L\���`}*Mk��\���k��O"H���Eڴe9�ndQGi�>���c즱��Ң���e��I$�o{���{ң��R_Cj�#��ܵ�V�6��	����2- W�k<���c�����g���Zd3ԑA�M�hWm�SX���n��D�6��-����l�ѥ�U,"�f,M�^��[+���8�1�&�M��e^e�/��=u�@��O�s5M�?�{gn��պ�k�u��Z|��u1�t��"
r� �G���偈�?rw�);�шE��X��{쥣j7�m�(~�H,=��j%_��XlxVHYEB    b631    1a00�=w��:�"�/��U�J.Õ��*�n��[-~Am午�����6��k�t71��2Ę,_g��2�N�v�J�Q���_K]�����d;����� &��r��wX��Nz��,
����|sQz��R������3a��S��q�;"X�'��5�ϝ,��.�
H��^���7{�s0h���N�Er����~:x÷��4peH�����ݖ��'ެ��mO���o�m�_��)�f�.-`�]�D��d�~2���6�`ˏ�?�����ֆ�]�q�x�v1��^	l��x��sC=g��Џ��2uU�8�g�I��f�e�V�U�͝�L���,Bt�c��E��P�Um4O�.G!��J�Q��}]�1z�1�ȟ���?�@�s�>%��Sb)�Z����%x�Abǆ�3����(�e�~�����4b�oZyە������&��t �D��8�-Eg�zkIi�ϲ������1b���)��0���k�qn���~���͛�ڔ�`��`�:��^-+'�'؈�` �dit���o#Ju�l�av<ޒ�9������D0�Sp.�cD��k�:aZC��	�z�F��w���K�d3�EԢ%'�#(�~�����/�e�����jn�6��@�3�e��_<B�ɟ�Ux���D�3ӧC2C
5�
g:w �o�(��{3J�n�Ƅ]ڽ�`��M3�:B9uŭIR瘏�z��Ei	�P�q��{��H� �͠�G_���kYCo�v��`�Æ�����I
�1��UsZ�v���pi���PG���0��:���i�#|��9��O�}F�f�P��������@&Ti���k�P���k��G��L�&⼬�imH{$@�l�:"�2G��@l�k��m�#S2@NAq-��^`�V�8»�#Z�`C�>ن�O(*T^��h-������/���'�i�혋����$-�#Ս@B���BT&�ϟJI	<w��gd�`���%�؍a���f/�s)nK�Xs5��V��
@k�֑v���UC`�}����Bz
2O��M����&�8�U*_�Ĭ�"�(�9MK�"?����k)��W�����e���}`�ƥ�pv���]m2�1ZW2]wD��Q��W��1\���]�^#��$6�k��jͪ�X�f�3�����6uT�qs�y�NY|�?$�♓�x+�O[�
�/�n�]�Q@/�EOZ�������`;�U=��I�|婮�4�n������쯯	�I�t�qp�D���S-�Ĭ��	Q�W����J�1�(�f|�QOڇ+������QmDִ���Z_^�e>����J��w�RA�|l�_��j��ܟԀ�5�}6Y�t�[�ߴ�y�-v�ùK3{#KD"T����"���la`}tnxh$׮��j	��~2�\W ~?7��f5���x�D)��Nd�o�O~�
b��C?Z�����E�+j�t�!�����n
$�a���p�hR��+r�O���B�gc:b��`���d�!�++��B�zS��g|Sb����/<�0
 �"�G�"��)���۬�V�8��B�� �,�a��awd�����UUޕ*���Nd��
(�ɓ���5�\Fq�}�sK�9�Y�S�_2��8�:Q/^w��p^�tB���4�W�n�q��� �"�ẉ}j��4�e��m����]C�o^-˗���7es�!$���:�+�Q],w�w����%mH3Y�``Ŷ�Һ��kQ*�U�.�9�x��`=�̳�/��/ ��u�S�l�/����6)����������	��8��]&�]�A���5���L1��y?,�v�3�e�+� ��TK��
� ������\�����d�C��\�bȎL>UC,�G;#� �8�ܹr�@l����q�Sv;}j#���x���9@66@R�9�aC3��M�4���*��#E����-�b}�	�OΉ���?�w.�ʕ�����4;X�܎d�޴) JZ�%��(��G���p�n���U�Ŗ�u?�p����G���	��5!6jdHGʛZyQ��Aѧ|^���{r@NB(@��?�݊��QH�C�U�"i���u��N�zQл���'80A6�#�5�v_ }1:���ݝզ��xS;��T퀠 V�!�z�g�+�=�JM�,2{.�K����m�/,�is�	Jx�]�_�=���@��GE�xG+��u�8Q�k ���Ļ%�
L�a�3 ��%[�]Tު�p-!����5�z�Ub��=��l���1�_�:V�!����3O�"��Z���2/o�b�\�٭�3��1�BQ����2�F��p�������`SOb���H���m���,f���� &�Q�`�6���\C&d�9k�B(o|��;����f�i2��@̙�G�/�-�z"����%('u���L%.m ꓁C��1�3�C��YM�@�����:̅e�G̾o�(+/ލts�HI�%T��}ة)�t�p�� u�/�b��B�rd��B���I����������_��	!m�Bܤ����B侣�{�����Qp�ćy5����=ؖ�+iKxt/��`N6}�}[�)�'�(����:��foL��w��,EZr�_-�&���#}�'�sՎ�@`��(��>iktR�x�8�pX�S���n�oOS�#��GO,��knϸ��{$Gh̰��6nPY~L�9�d)^��2�o�|?�ͤ7����ã�,ܙ-a� 3�����E�O�a �8��$)N�ms	�TjG|�����5����ROZ�����[��M��D*.�xt`~���>	}Ā�Âu'Z:�E�$ް� �n�T��a��3=���V3$KJ�x��֠�+!��iOc�;�*g�e������`J�RS����0�H
+���Q�[Y�Ͻ�ˀ���&�ې�L�� >��4�����!ئ��:A����ccaQ�o��<����\����.�|�O��1y�gB��������W?d5T\(�Ɏ�����d^� �'O,,��������V�zP'gCu��WE�lt2�GC	b��#H3�Ϝ���Q�O��娣�.�%q��rhۺC�5}m 1�,5��/a@��6�
��{~�WӢpdu��rC�p<9Sj�ܦ�e����U�-V\+8��m����P 7-Յ��l��p��j��d��)�9@ϳ��IZ��!� �5����+�Z-��?��<M5R�eH��y������y�Ƕ�D|W�5��Ut<�N��tг�����k ��pb;�/�YҸ�椉y\_�/D�h$Z�Ԕ�L)�G�;��p'��P�"��}~��{f�yvh8R�LH��^����f�"��0dF~0�5ǵ��[�!�H�`C$��V�)�6�>�r�����":}���B����sYw^���'��"\���dìS���ŔZ������F�əb�iz�Zj����$���+_���ۣE�����Hѳ^*�84)��pڗf��Cw�ʁ	 D��}ڕ��I�JދSD�I�&�Haʄ3�@C���b�c�����_>;}_s����K8�˯��r0�.�+��}�&�3����o�ՙ��)p'�$�K��T�me;�D�hq�O�sr�8�&.QQ@o{�x=i�Ѝس��\X�V��M7��Xժg�^�?0�Ms��['���KT ��y�C�7�N���j��0˝e7����M/�ܵ���꼠q��QYK����H� �c��o�f���-�#��>���G����*����@:{�������׿��� ��G�E��~�5hfK�������4� �P���B���~J#�gXV����jA�5v������E����[�2����IDx���<�I�j�ߚ�� $ړ����afVb��/�g�W���8�9�Ί�槸�'&%Ί�j�@������[�|$.V���c�H����^1����%�"+�il��%��Z�v�R��h[�3��,<lRI��p�<4R�Ƭ�%p��2t�K�7<}}�vl�����JD�c�Ae�}�0�s<L���ܴx���:��>��P&�IpI�o;�7a�������X�b56�PϪ�����]d����t���V���ԓ�������N&�C\�����u�q���n��qi�a�������TA�eU�LΠ�lD��'#".�#B�uN�9)1.��kG$�u��f�D��a�%i�r8*�m[Nv�&<�;5����F�C�زBec8���ةNk&�?�8�v&@��/�� Ջnb?�$WQu�{C��ws.��Wk�-T}u7A5!��K
Ĕ���f���k��ht�m�l�8c;E�Xj1���\_����Ž��OoK2�O��@��z
�J��vp��<��ʅ[m�RXܐ����<����
��:�l.��.�"2��Ё�H~;�j��/(:�b�}��Py����+��8n�.��*6I��_j�A,tqN��'�Gg ��|���#[�A��3���i<sV}Hk�FB9�y�������)�_�+�0�����
�4F�$�A��M�빚��x��#vRuU�k%g)ߐ������iq=v��~�d����?�E��z����O�׷����K?4M���yܚ����>�d����"!!���Sē�c���`�r��v�'�&�o�)'�JB�i�볔������~�����و/Tu�������M]sq���/@�U�<�f[8�-i�/��9?�jZ@�]��]�P�GQ�'*j�-�Ÿ�aƿ�	��a��,�ø�Z���t%�Z蟂��@���@*O�����GN$cV��	���
l>�O6���t���?u/0��M4�i{�-|�\��?h�jJP���������sw�o?`~�I-#���9P� >jK��5�vr���3���5ݔ��`:��`�.N[���2��_�����GY:�=��+�I��T�r4��^����[�#��j��{�^-�Z�_=Y;�_娼k��y0ۻS�િ�L���^8�50H�uz�3|�r�U��-�|�^dV�3���ae�>Y��]���D?�Uvt����d�K��O����5c�a���d�J ���Z�C>��QȨ4n�s�p ��ytG��:����x�0�av�X�rL$b�U���&O����r��)��j���:��q[(:�2K9�f�~N���H+o)_nZw_J�`�7���9A��n�������{��w�X�e�>�-�8c�o7jr {/���Z������6;�glw�%�r+�X��Wi"K;�ܩ%��t	Q0ϖ���}��ɯ�m"���3e^�V?/�������#"w�����mꮱɈ�������I:l�		� A��N�}��F�<4�n�֌��@y�,?ZQ��?f�^ �oCtA�f1貺�e�	��t������XZ��g������zj;x���(��J��;1u^!�4�,m����R>mmL�;�6���%c��V>�0\��B�{�Ms� %����WG�%';������Ϩ������-?mu^�o����5���7cl^\)�G娪Z�K�U*�,��H��?�fJ���f��8ܻ���d-�;_�EO�9EG��s�Gy���]4��d���4���@�9"tJ��4�,��Lmc+��N�:0��T�
V�^���xB�*�R{��?m��cO��.�:���:D�4T��b���XDx$\�����w���eP��e���M_V�:�t���1�;&�Ͻ*VS58�֡�n���-hP��]�S��,A�t8)� ء���+psӆ��:��7}j�% e<<�>Nߖ>$�vO���Cc0^��wp-�;����������޲�OK�����GҪ��0�Y��>����$�&gS����H��S1���حC��1R%�|*����EnRp����ḡ����1���`��]��vD1,/�zA�@��#�n�6́��ڞB���7�����a�T��?f��cM���WÞ࿊hZox?l�>s��\�V�X�<!7��]H�<��U)��QN��͒>Sa�(�V��v}��i�o�b&VYy����Y�,Km�{uNi�r�<���TB���kUT�܈�qj�K#��g�{�D���%��#��XE��O��e���{R'���ǩp�w ��9��yu�{׷���t}P(풢��!�L���)'�\O�Y�����������I���oU.C����U���Sw���Q��@�����1�)q�z����Ӡ�Xn�U�;���\�]�!�y�Ƿ�7~���c�jR�#*��:'ړ���)�	�U~GĜ"����C�j6����D����Ƣ�4�~ބ�}6 m �<���'Wh����i�EY���͆�S��2'��0��.\P�nb�¹�B�Ί�(M�:!顗�ú�jy@���K(��L�T\?L�G�?=���)�rw�?�U����&� Vâ8�,���wg�X��A'}����ı��Ȧ�����3�wߨ%�<�Bp�5�#@%2�