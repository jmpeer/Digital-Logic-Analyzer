XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[|(UPN3���F�������G�
�7�K���'l�L�� �m^j����0[}��0+��E�ذ�����.Ƴ�q��*� F}��2� �u��A�.<���'8i?%��P���mgIbI��>/뻅>�u���!mC{̛�$���&i�61��4�@%>L��5�4���Lr��svnq�Ԍ�!�z;n1�\":/<��ns@��@����;Aot�˕��R���r�U�	������t/���H�6�NQB~��.���5��ڲ<}H������hQrT��)6�e�.���C~���`�$�HBGޗ����Ӻ�;�pҚ3|#l#�}&�o҂%u0DZXgl.+�?��eiU��S5��$٫�ӡV5�dڠ�H�������鯍�y�34W��vs����]�U�4�BG{�1ox���pJ��  vL�E֣�g�͐�$���vG��X:`I�|�v����6�E~��a��=����X�Ѕ���m*�2�.�� ��v��Y��V��}�-�M�f�{N|�=���"Yul�}�W�h��x3qg@���W��pm;U��޼N�g�4���ן<���#�������{s�� ݹm�Dk[�ׂ�Їi��_�;c�w��7�c5m�t 7d��uՑ����J�$� ����#�=y���Ç�<�
1�ڲ��m���P���KB��q�ɣ-�
���ʲz�{k{�M����lj�i�h7�4�����u���ŷ��>�ccH���:�B��AXlxVHYEB    fa00    1ca0���.�\b-�H"����ڧ���~UE� ����������"��Ƨ����q�,[�g=�IقЈ���]\=������:{�(�-����'�@p:(:��e�y`F��Ҩ���fn��O\~��Z2�����n��|�����}�������䡬���2{�u0�F�'�ޡ�x� A ��!��>�k�t�.��z��ᣲ�X� >(���b@G߰�
��BY����W�en��S?!"��rIsT�#ڟNd�3���ꗈҽ���O\��Y�8j��E>���RQ:BU�r� �5:\��j�_�B.?|^=��� c�J],�c|/f^�KAOyr��#���6EnY�e�S&��g�f�\M�2m���C}5�_�:Ve�L�d���F��\ii1fG�)����� ���"[<1\��7�w�>��mt`�M%�<�9	/��� �@Xm_��9'��\o��1�/���^7��0q�7 9uv���k�٬��}�7*�;�tDF����/hVT�W��)�I$
��?� = 1mgo|J�o��>�:��DÇ: m���G���!�J{9��;c�f#���K]}�ݫ}��9c�u��9	��p�t� �dDpD�J��z��A����Vr0��ZD,��I)�C��Szb�Q�{R���;a�`
c8�-�F�8d�P��������r�B�@	��-p�����m���!Y���	���o��k�:���(��7��Q
�k��U�+�������H�'�?�cM%?UJ�a�����o�D5֦�4�~�v=��{�?���fρ4TF"�������Z�y��8~#qf�Ӧ��� /�N؍'�k���=�G���
|��,r'd�brZ��h�Q�"��y�.����֒.m�#K]�5�0�M�BV���DJƩ�sR@Z�
fX��(�O#�.���+�61(�|�xÉ�����Ɂ{����y(�c�rzN�1��D��^B������ƀ��1�D
M�$S����a�#Ԡ��i̿fc;�!�ی3)~�m���)t�:�s���זV��E�!ۆ b�v������gƇj��_�L0 ���v!<�_��63�}��'>T�/TI�܈�~ϒy�3�N�3�.���I�K�*�"̠<��U��|����\��}�`��}�DL3fg1$(��{�|x�`��_	LM��̚;���ɢ����r0���@�-xAT�oN����8u���[�Y��\�1h!�K>\����W y/��JZ�q����4���f�x/�^��:!0)�2	F���j�E"��|YC8y��R�U�W�K����'ʸ�1��{'���B�I�I� ���F�.y*ϐ��❀V�v>���}���`�ɘ/�$��S��-$ �W�!B�ݾ'Fi�8B��15OI�T�D��c��]Nܮ���F�b�Kԇ���ni-38k,�9���R�t3ZR" �=t��Z.��o����}j�\U&�V�۶t�N����oW��٭܉�bd|���@��k�u��B�J���&A�I�u��6�A$g�Q=�ܥP���*�s�>|���:����R$��W(�)+ ��(�� 7�:�lw^�ܐR*wq2�n�)u�ꪟ5��Oo5��,��G�O�n�p�i�g\��;��r�y՗#�u�#�3����7�7�i�!V�{2+�NU��T�_-s�E��Y�):����=�i0@Qۍ�)��o��Ǟ^��df�\e�o�--dڗ�u�0 �̗���F*�B�t��<K>!(��K��RE��@��׼WA�*����-��]���\��>�������%���*��6*w���M�Fz������T�vM,�u��*���
Z���Uaq7+GＮ�}��ު�<2��|1�B���Dk�o�.j�_/���yI��	��N��*Gj��W�tT����r�\(Wc���4a%o�����s���"�θ�\�bs��ѐ-���X�t��}3���T�}�\�k��K�%�N��SϏ��卾E�����hI�2c�]�U��{�m��'=�������T��0�Δ��/.�S�nM,3����"נ�;�e�g��MU�9N@��j�-��o�����8�c��B:�C5�3�
�!@�u1�R� w����P��Խ <|g@�⽣{�E���#rD���^y#�k4���iX���YE�(qXi��Cg�2��u�n�w1��-�Ȁ;�vt��B�'R�(?@�ᙃ�����uS����Sӷ?��8m9�r�_��!��X�o�/qV0j)��BS�s�^�ߣ$l-����Z_����Ȑ�bk��+��=4��e�`�߅x���T��H�Ӈ])��E*��a�%Uy���$�|*x=�(F�K�$Q���C������	��,9M}og��I�/���W|�~����?���>�J\����u#j����W���.6�`�k|s-{�c���qL5�1��0EE:���ɞ�,~�`|�;��B'�'\�j����OL�,K���l���°�"3������Y���Q&�6a�`I>�7(��N���T�Ɛ�c��Y�2[�+�ۧ�C�[�ש������{�	ϰ��E̡Ժ2��&[�Av�$H>�%�����bA���@� �ogG�����[S� dA������jZ@Pa-�S��VZ�^ۥ�lV�^�O�w�ʽ��O�W�3~_*�7	'6�k��!����(���R�w�WR�P��S��R�m1_�{���k'�ѵ�~6�Y0sʮ�a�1|G��|Q9�
�W�yA�rh��jgVU�f�\�M
r�K�3��� ���MUwr�?^o1�,
,8֟p��#�&J:�߇ƿP"ǝUi'mO+Mx�F_O$��������Q�����Q�0FAB�E�Έ�5}[�
rw�9L�e���� -?R������'Q&�G���;���.��m�@7Ϸ>5��]je��Y��8�Q9�b�"���X+�i��J;i��!L(�G��i׫E���Iճ�d�.�Gxܶ������߭�����[M�"�ٯo�1&�qws�i�t�G$�\Z��M���s�B2Ϭ5��h!�B|x��n�B�}�~|�#�ȶr��ט��9V����d�c�j `H/W~ᆛ���ձZ���'8o����^ Q��G��lP&p��qu�;����Î���y�iJ���եVC�|bՙ	X�_��B��t�fQ�@J��?	���.*���&���+F��i�*�7���y���q���0b�2���ؔG�Լ����3��ẽ��&Hc�=՘>�d����;;�"�ms�Lr�a'�U<�����	�M'a��%�Jʕg�O2,���7/IB%��0��h,�blvvaY<�,�]q�g���^|�4ڛ��K��s�ZϨ�I���X�N.�]p�С��ct��;"(�����1�K爊-P�C:��W6�磪
�4�8��$֣��Mإ1�P��j�s��݋����b����ꬦ�uS���aF�%}�Ok�"�"�F�B�s:p�QA�;�[4q���Ou�u�,'�
]�Qx�La��2�0��ƀ���sNz%�Ŋ�3I�_'�i��;,�B�_z��T�{�Ծw��<v6j���J��7���@�6D-����z�A���(A��m�Q�^\��:׀��/�Ӌ�?������۷.!Qd���#�W���r.g]�'�Gea"c�;ş9F/��ɍ�S�̼P)��:^a��P�Y[(���l$�����5�WK�b��:k/4�ʮu�cxݬ�&I�(��MB�J� ���v�����ˍBpt&��rYf�y",Bm<!�x�L���_��}����B��<R��DДX��������ˡ��z���\ϳ��YFN0��re����;��'��p�E�|�1�c�^z������?Db��g����Cօ*�C CSe�+��i�fpSvy0<C�c-w��;�4qq�)�&CY�+��au��!W� v�L;��EY:rցϒiY�}�?tpl��ꎔ��M�,���3n�|*Bf��6'n�׾�x�O����wi}��y��j�?�����I�%�<E̻��tp�����W��n��Wd�+��3-bL�����EV�l�����a�?[�� 3x{ ���6�l������>�I�gqq���ҁ8t$CČ�C��D^y��sU�+��]�@U*��,1����z��p�y���F�|E���	��-	Dt.<ضQj u�%���!苬>�Z?��Lf���|�#��\$JHK�6�UJ�C��i���S�z��C2�RD؟:��aCㆍ�j5�vnO��)8� E�CL��}����D���~^]<��4F�%��^N�zy�E���YX��+���;�@�+��-�?�v=�X!���"fJ�w(�����1��p�A����J*pGEm��><����^���r���yt��7/5�<�v����_W=,ޞwkn�r<���Pҍ�j����I`�j-����˪j
���QI�sJ�����35����(�m��f `����D�pS�oܹ2D�� ,�
V����)��Q�c`z��k����ry�k
�,�+1�Φ�-���*���>76?��qaO���v�wL�r[J��G�h�Mq�(ĺؾ�5�mcTv����c|�6BU�ɹI):hd=C�dq{�6k���8���d+rX��oXE�+��ʏ-�E���t�#��f�w�e�H"��5�-���?��2>)lC����Fv�{1X�Ak��EYH+��Bv��x���%���4F8ޛ��O(���=��s��<\���*A�	p����ЇTe�j��[��E�}	�:l���C��4��9�K��1V���j��}~�����*�J���G���-�DZc)V�L��<�@[5��!��4�0�b�-�x8u��5������+6��E	�,_�����o�)�7P��E!�l�+�F�������Q����� {��3�C�
˙v���	地�W���PPSn�&Å��I�M����@���(Ȉ��!�G{j��ʀ�e]B@�+лth�O���,�9�k��c
�ҙ�B�G��1�=�mQ����0�]O̞uk.B;�1����-��?k�jp:�L�s��w�>y��J3��F'f&X��zKLJ��)h�)t+U��B{�!*؅ڄ�Y���y���1�uz��I+��mu2-�v����"GQ}ʬ�V��zH&��ԙ�`��qM��\^��;^�_�>f��g�k/�	�Ju�����.�j��P"K[:,��SBe9l��)6��&������)a���6��r��$�S��m"�l�-��{L���,D�R��V��ǈ^_�Z���u߅ ��x\Q@go��c�9�����]R�8Z�@ ¯{�T�I;�!P���b��Z\������1�c{�j)B3*��X!�hl]�wα
��\tW�B,?���N݆����GZ�>�=����`IU!v��
���ы2˴��3wơU���Ny��'j9���gr�-ɜW�S�����Ο�����l�b�T۱���-��wC��'�@0�B�-�Ì���>sN	���P���;�p�Ń�w�����4u���=>#��$-��k�{w�B����d��带�F0W��ִ!��i�����NΦV���u?S�p�l+-� �8���bO�V��S�)�z��}]��$���+:�G����;?~�R�� ��Le`�˜v� �P��]��_�_���Xg�a�K����H2ǘQ���[�~�jM�%g.�ѡ��Q"R�з6��\�W���S�7�Z� %�xN�5�Z���:��]>����S!�#�����:���ߞ������j�.y����� ���R}'����4Hӕ��*�\ML$�u2XHv� ���8a�����bS����؜P7�š;�L�p�H�<MW/ 0m�#�7V�fTZ��JK=u׍ѫWź������^k_�u,s��
;eKB.����q�Q]\|��y�;���t���9�W�ڥ��\�y��+����8əNP���<�@0�"���c<��Ꮄ�����G���?/��]��o(g'��/�u�`�~_��ӠJ��
p8��}�ܝ3{�� �����D��ă�a�QV�#��f��Q�2�,ҽ��ķO����2��ѩ�jE҇���l��@�ۅ�=R�:���&���hgT`$X���:�
��c�9L��	X"�N�|(�{�|�Pf}�0���r�N�-�Y��/A�V6i>��'���YA�/;=Ij�tC,���H�4�͟�/_"��;##9`q��FߎBa=,q���JQ�:�7�W�+"��f���9i���}O_er2�U<2�j;o1��x����`Ue>6�s\y���x�JU`f)�N���@���&2�J3:��}.Nm��	�pH�KVӁr3<�!_��u_�Lvv[[�蟬�6 ���o$AFy̱(#���҅�ؚ�^�	"���yM�2��	ke�E���� ��xUU&4�n���%�J0d�� �r���.����?������ޒ�~0�$Iyџ�H�ؤX�����x�0�R�
xp���7nm�y��'J:��W1���<�6Q=d��L�Z+���/;�ή���t�Vk6k�a/�Gh��;#]b�j�)d�9	XF�kCh�1�?hTY��u�m�Ay|p��~�������o���[�p���,�vt�ha��7Q�d�K,�������&[id�2�̫��{::L�� ��J�"8i��H)Q�"q����0��n#����0���P�5TZ-�3�$���P�Q�X�X�3E�OYv�����s�����7�i��g��Q1Q(ÿ2��VS�}|�g��QQ7<:O����)�8�L�Vʢ�h!&�9ej]eR��޶&Փ�����J�lBꡖ�3����3�a6Ĵ*�G晼��#|�s'�n�<kN�lt�!��.
*�4�sÐ<���fndQ{V��ap�V4�=��������Ixi}�)�lV�����>��~6DX�'�_���Jesi�ڝQ{��\O<;C �e��%��f<���]E�(�� �T�-�}��dj; [f49�^n|;:)���W0AdT��L�<���;-����6�W�-XlxVHYEB    fa00     cf0��4`�����MJQ0n��8:B��l����l^����JtpiG儿f8�9m��,Y���7�0��Z:�N�(��a��
�D��vm�b�����m��M�3�Q����2���.l.�m�bj�tt/.M������

ܟ�[F�]�;��y�ϥV�v=��#��/(z�)O�h�Q���ّ���R)� ��n��;�T�}�'B$1E�*�^;"K]3����$P�~+�D��D��e�*��K�P 0ן"�9E�AS���~��5O��P�)��� >�lO)bؠ���Jo�l"����]b��s��<�?;��~�����52t�[�ё�D=ͻ_f�gH�
�T� �~�?!z�K��hl��8JSn�7"D�r����=Ӣ��B�푏c�X?g��>��=- 4�/�*b/AGV0��=g�cIND*Zg*�F	�'�$Mr�!�Kr�{:$.aXp�ϊ��̪ן~>�D�ߺȱG	T�V�{����Ve]�*���-�&�d��_0�b̻�/��;Q�c�T�Ĉ�Q�'���R-R6~����}C�a���9�.L}���E�'c�#R/ Wv��J!�G���*��`�Q�+~�u:�5.����$���n�*�[��H�|�>�}䴆�0�E(�.�e�-��~زo�>"�,��������$aJ#?�[�M�x�W�����*B!KZ�51:M �o���}t����ع��
e��h,�Ij7������X'�%��呤J��!�T�w�x.����M������$��_.����?8b��^�k]��^�*Β�|�>�Ka�gp�Dt��+`��.�lp�b�.PR%q�+j�3�ǈA߱-A+F�"�m�hE7 1�sDڐq��ɽE[�Tf�9)'�~$�hb�ľ	v�`�	�zw�"� ��j^^�󇱀P�~8�Z���$���	
����Q�nsnÇ�m���;��5M�J��>����`��$� �i��gM2����Yaǝ�B��@}񣢎��s��ϓ����~��6���;���|id���1���i�S^��
 4c'��ďQ�g02ZM�NY6�����n���� I��]u��h�t�Y<ZM�,H[3��OX�:6�:+Y@{�y���1�k(|8�9�$tݽ��I�hwC_o(Ch�Tu��@���� ��~c���S����#�x�ɘ��ʣ@�h�{��c��0��2����$��L/}�:��V�je�Db:+��<4-u��wE����w6F)�rtv���n����i�a�b3�<kj��>U�>.�b���T�c��gr�a���Xƚ�B����Y^gyNIb��=s�1�����[²����Ah;��S�1�5�5�A�j�\R���o��$�Y�W��B(וڭc|Q[Ԯ��"�>H���.��ܦ���˟����=B׉c9/�ZW��;$ڠ�bo�PZK����0���B^,�
Rt�ֿL~�Ey���'ꉫ��b��ד�.~����(��T�#��)�[-�T�>0[�����+$���l���o��� \�\�=nU3�l:�k���~�� �w��}6o���.������%�T�wQ�i>z��|��}6���j_��u������C�����~�Rf������������mӐ��$1pv8��]��/6��{,�2�����n�%��1��\�u��/�(���{��M��R��$�(�m+��_��r�����£N���ɛ��+ɖ.�A��Kϙ��:H��C;�������.=�3���8-��Ory�k���u�i�=� ��b�{5zv�%L��rq�|�q�y�&W��k%|	�/���>���S��xU��:�
ǧ��{�I��� �-(^��>���حJ�v?�vP�󃸚B�o�� 	�N𫩛p�!�Xc�h�x��������5��I�@R��aB�73��]Q@��%������7:��4�Rtg̞�T�"��t�a�IyI���y�/��4K�.b���&)Kj��N�O��]#d$2���� ��2�lH���+�m�n�0><\�P�U�g?�����ϒ+�@�̓�MDE�����)$�S����ݐC�sI*D�e�[]��x��Vl"ꊂW�6�oٚ�x�O�U��މ�<Jܩ���ަ��ۅ��L�:=ѰR��>k�U~��>��3��S�RRf[�������!}���
!`.g�q����J����j��@.U!�b߂tу�h��K�K��O�Z(���ó�	.y� " �:Wl�v��Y�[�*�3c>]d ����֔|y6ŢN�Ÿ�I�1�;����W��V�������2{��[����2�}���U��|��^k�=TS�̕��	��]��uܮ����p��]mZc[m�����y����XqqOi���#~w�u6�)���4��SO����+`��&o
P8G£ﶛ��{�ײֵ����R�IZ��s�ۇ'`�J�ߊ���f^�N�K���L��}��I��l�<Y�A��p�����V(~�,����+K�^�X�2�/��0�ܗ%������[.���ܖ�H�G3i�C�q����/����c�̾//��8i���1k�ۘS���A,S�"�Bw�� �V;R�M8��f(K譡�qgf!��,:���k�����F�l�h�H^�;��/��7��Hp3
����ľ����F�[������̦O������۳h�F���WH��=���*��[��
��)71;����6S�+�V����(�8~��7�A�Μ7��r�h�|��Σ�E��bF�� ��0&�~��є ����ŝ"@�U�b8�4?��V'�K� �R�j#����+�y�ľ�W�A%D�X��d�wGa�'њ���O�K��@F-��n=Z�\U�Sr�a�Y$BsӸW�;*sU�g>�1-��\�+��7��E�3nF:�MUAy�!\(c�j�� �3��F�ݑ��2X �˗8���a����o'�a?F�w���a���Gy�\����ae�r��hE��L�X��> ϰ�A��=ǜQ\���a�E#8��|��8))^��B���5�r�h*���`.[`��9d�zq|T�����'�.����C`I5���叏�3�z"���CU��!.	_��Й��ܬ��H�s����t|��/�wU�t����"{z�\�7U������[uO1�2�DL�ejC�S����#`nr��20�� ?9�.���G���:n�pSL��­G�&�����a�IXlxVHYEB    3981     4d0��ŧ��3�0,� ���9���{h�y �n'O��d�
>�
�[�{��|r�D�T�X���׸�]��Bn�bߜ�J)��:2�kê����r��s�TQuԋ�Kei��>�v��q��
�a#��N�a:"j&QL����׺��(<n��`�.�"p���oU��c���x�9�u�g�-��Z���,H��яȓ=&�,]��qҒ�wCܟ�G�_c���E�ύ�C�O�&I�1N����eՏ���b�l��{ɐ�t���a�"`�ۻ-# ����ؓ��D�\�����^�Q�����pBj�^"4��s0D[F�_e��-l�pя�O�-�Sl��li߲�i��nHk��$�w�6�Vj������BbB��$V�@�ci�-�>bY�I���p��d���';�en��B���/e)�Hq���-_%W%�4���$��Ҭ.�[�sՓU���a���8O�.�E��a"E����e��oW2�Pp�L8���w�� ���c�H[�R���M(��CR"��-J��K��Ð@f+�w��mʧ�g�j�͕�WR�3�Xc�'�v��GG�o�P����*\�b�(�"#ɇ#9�� !���k�P&�L9�T�cD��"\�r��w�*����x��Z�V�rQE�����	9)tޛ�bl!��,t�Fv�dD�H��b�`ןvVY�Q�)Q��ɵc����"_�+;p��S� �HJ�%�h��L2�@]�I�}����͢��(4���*�ڰ�nb,b�b�ͅ�u�U����rR4���Q+"&��}�Ӥ��K���}�j����ay�r]�(�D��	fH��y���-��t������j&=x�:',�h=S�|x�pN�w~���.���QzN����Al�
ޱn����L�o7zb�Ӫo8\��n�p#]i�i�󴍾*[�ASV�Z@�z~7�g��v�'�1`�q��V�<�t
��J��Z��}`���"֊�xԡ\�>���w	�F>�W�aQ�v��� Ƨ�����d����𺞬s�
�;����2��T�1Ϭj�׺,G w1_$ݐ�MM+mcQ��D6�,�md�j��?Q��w6"7�B	��	��y6/����ʕ~�}r�И��NB��j�!��A�?^���	������:8`ָ��0�0�J��������ȹ� s�� ���%��Ǐ(p>�^�q�+J��x۰O��