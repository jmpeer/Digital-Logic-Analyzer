XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���0���\���L��.��]Ҩ�#�m�1^iGʙy�������
�/���kK��fu�}3�V�\ ^+���S����)�����{.�~*�E,�+�~H����$S��W��'F�ǆLXѳ�"�������+,� ����İ���n�������u�{����r��~Y#\�)Gse'���W^T��ռ��pץ���0���f�i7�ymw7�G,>n.�`�0s{s��'&���|cQ�HBL����+[�C�q�U�5�~�ݖ�Z^�W��h�� ��Mv����LI$a'�E����S�fF&
��T�յi���e��@��y4?C�Y�W�@7г8�K�z�eu�-�{:���s=_I��U���-C ��N�h���J�Pj���*�+��5a����洕���xA@2)��� n� %��;2Zl���H��u��`Mou>�q���y�%�-]�x5�>��X�n�W��kn�fRd�t����%@�|&*��G�$����'C%_i��b�Ɠ -қ<�wb�� "�;�~^�aI�t{'|�U/"m~�g�r5��_�J#3쉠�V~��ֶ~݃��n�3?mz�m������3�mN�L
���R����`����I(�����Ζ;,��x���˓ҟoAZ�=H����"v�B��}�"�))�gk����X�@6ȱtw�MY�E�N��l���u��1�E;��XS��4-�?q>Cz�H��~�>{mդm��C՛��}<�n�@b�XlxVHYEB    fa00    2020K�} ="J�<�KʛY^r��ä,�p�2���5T���W��RY�Q����5G��C��Fn>�<0�R�=<�DT+��Hu89�sc��<=���,���o���h8���}���ٜuMe������۽�Y�	�A�*�l���p_�%$c&���8h���E�F���8�H����%���ɿ�۵(_�k��w��0�țE=���2���|$�W�kA%��
t0A�2}XS�#>�mVYK	����fTX�iav��]7�{pJcs���0�Dθ�><�xN����A�.�b<TeE��AQ��z|������Tr�)�<��n�������γ��v}���F��2#(�sqOM׳+o.Dz��@����W��n�`�K`A�<����	���U7�خY�����Ӵڗ�1�;Ӿ��&��O�ַ�@�<�g*R$9��5��9�)��P�1�!�Qo�`+ֈH���\2�<)@"G���vY����wo�}f�1�3ˤB��	��Fħ��`�����pyHD�f^�ߚ�+�r���̕�Q������vX-�/�/rj��,W�ְ������8PM�]��?\O	�	/뱘��T��=�Y���_B�� ���#"���O��ZVؗ<��4x�D�`^:.�GU�4A��;EL7���|����cm�	RF��]����3�N/�S;ǟ,%q#(�!	���+�J���X�i��+���:R��D�Efdfr��/��Y� �C-���@E��L�Y��}6�sN�h:[�>1�Z�z���C�O��:�-�0��FQ=��|�F���؛�=@��4��˩h⚙� �.}#w މ�B�:d��rx�g�p��T�3*���	GM#�)��JlU]�|<{�n��̌Y.�d4u���-�XC@c��`��adOdvy���_nR���4S��>��g�&S8���(@xh%'��M���\R��GFH+�`��J��9`K�N�Ѯ�(�/<��kƔV�%�ca���~n�K����������q"B�dW0�>V���'7���s��"��j�X�?�r���i��򊆱�K�����ʵJ�!�B���$R�݁�4m��5y�>�JKp�s8�<�Z��Z��5���,(���^_�P�����"�ae���Bi�I��[`��[ %Rs!�@upC�y�V�oVz�UQx�Q�F���C��a������Qq=�-q�+xaU�^���<i�
�ʹ{tg�s"��^N�]��=�[��6�wi��4 +�FB���e�}`�:����6"����=?�<��޷"�KD`��K�2����2�ʷ��wK�<�B�	��v
�c	��)Jr5�u[Q���qX4��ݥ��ڋ�[
 SD��Oڻz�ߏ�gl���X��~\Z$��D��̐��dvg&�Z�~�Ja=4�����;��:�����z�!il,�T��ֹ]*��JU����-�BrbM~�w+� ��/�21��S����gŖ¦����.Y�eh�c���a�Bi7�0�z	2�G_�zۗ  qc,k��y�R8���i�ډ/���t���R��eW�.��Q�̘��Ժy'��?�P�����Z��E�ǈ�;��̰��&�c-��o|�C>��������rL�A���2���X�l�p��^<����q��n0Y�Z��C?uv�e�5*������>�If��h��-��Qڑ�s�^w#�L-.�B�g<S��T�PB|�ih�'�j��$���L@h��C��*�#��je�a��2�0@( ��@s�lSK �q��g�:+?����A��4c0��7��'�b�i���qdSV�'�T���6��p�*ѬX ��țR��M=�ޞձw��1�v�!>\u/Ux},�=?����͇�:��#�@ߺ�A0ps]ϸ�>ClK�lR����@K�ؠ��i6Dɗ�Q(������ы��8�d�<��0��HJ�*��1��x�D<��Dɛ�
ux�9BH@Fj�ZZ�^O�����$43��ȧ�[���f����r.����ރL��n�uᴬƿ�)��9���P�z�Y��̠]�3�m���z�o��tP�~�h�o�{.�� n�v���\�ܐkh�$��Ei���k*K/B�-3o]��6�Fg��xj�,+�tN]����~�I��C�u]�/���Ɋ�cz���gc._z�p�>y�@�=p�!vM/�ΐ��`�� ��6?lk��CX�2��f0�|�k��Ě����ʲ��	��T.D\V��z	1���8�������htJb!>��r��p��z�� "W[vc6�vP�� +���ڊ�n��fʔ֭��ʯ5"������`;�VIh�fR��I�<���<��� ~ϴh}e=C��f1�	�#���|��V�C�ϝ�w�.u�AM��pp��R���!.~�U�nr"w���u����׌�݉��၍�rp$KXa!�%z+�P;�Ӯ�+S;+����>���"�)�>��"x����������x���D��W��İ�H|!S��#%A�z�>9<���ŕ����L.�,^Hg�>ԝ�7�\�r{SPQCC,�4�*��[U��������}���� �
dy�d w5���a�H˒�4��Up�$e5A	|�6H����@�|:c�.v$vr���"s�N�ޒhW�U��XJ��{$ɶ5쮺��]�Yb�>65��5q5\�W�mR&���H�����y��
��~O/�a��:��b��V��0o��c�G5�y���(�Q�G���t�:���;�Y��GKG ݸGq{�i��:ƭ��h����zd�6pC��W*�d���C���N/��
��| �2V��9 p�!:�?���c�r�V���M�!�[��O��T��TC0�C��ϸ��ϔj8�C:�~�]6�x�E�aO�E���ez'����+YT���� ��c�i�o
t�y����]�Y�F%�w�S��sC�f�l����5Bq�"7�-G5aw�!��7@��@p�CO�˱�eg�(��,gTh�:0�e*TO@�S�=�������Z��j��*��i�m7B�����l'���mL:}���˝��S��r4�T�w qk���8R�nB�����]G�/Z^_�9�$}N�9�S8ɖ��k���C��S�'Q���l���/g��滇$���d]��)��_�ݻ:|����ء�\��8w�\�IE2�7$��%�f�����R��"���X5���+p�ڧ��,ȓ���	i"uٴ�\�7��C���w������� g��-�@�"�ڮ��0Fp����LH.���/��E<�1�E��0SЅ��Cc�~�\{<���1�a'�����bx�ǋ�I�+���&��6"44�`�����p��L׃{i�����ע�!��L��B?�}�7ޝ�ۓ_,��6%p_�Bt���6�أ��܋d�Z��l�(��&��8/�G�H�`��8��u�I�֭�̈́�O���AMНam#�r�����UQ(�M �����  tO��� mB:�^��ZP�"�w#<�0f���c�At�b��z�⚯C�:z�����KeI�s!*Bĭ�R*�]]u��g�kօL�#�L�a0�������Y��$��m���KK��;'���� ����
 �;����lm����o�޺ �ߟY\��L7=����G�7��Է�%_��A�W��"b=״�R==�G�����
*i8p�*h�Oj�x�cD�~趉�?3��H:'��{�U���JN��[8��P�7�͒V*V��I��o����p
-%q��St��t���O�XM�x;�ny�����X}4�=U}�����\��CU5�N�9Z����P�Nk��4����z�)�$�Y��p�?[���~6�1�@;e�0*�"��xr��*�>��1`@�϶��bb�f��,d�����a�����VVVg�
��̱���W��A��wu@�y[��7:x�ܺĬ
�`��eaw�y@#,�N�B��<K�c��8�2��L������ih%�����cC�6�1�W�b�jήr����)oqs�R|OӞ݅z��4��0�����L���U:��ú8�/����"<"A�2��2Ƃ��������Er��ߒ��n_ƿ�-�ޜ�C(����,�
$%��by��ՔSaF0�a<+����Vf�|��-�N�S`V��-��J@mӮ_uQHh9���g�	$F=:�����Ӵ(��VbeF�����8��������D��`��4��i�Iy	��D�b0���u�F"2ՃN�TZ�Y5#����.N��Ka�n5��Ѐ���WNPv�O�_��W;��{C��L�B^�����J��D�_3d��f<�q��"ő�D�_�5��1t[�b��k��(��=��>9L�C��!�Q�$9����|
�n�4j#������k\���g�VfPF:� S�H��߽�����kG��d��1���Ǜ�"+*D���/�v��?&g���{��*гHۋM;)�lMo�xx�|j�8A�R��)��|��~G�>Y�}��1^�J.��W��
�L�Qn��HHW��ϼ;�k!/<�)x�#��L'ϥ��� (�� �C�t�'��d-�I�m�|�6WQ�S��9A�x{�����z\���v��e�x�	��/!��P�a]iٳ&y�=�̯]˂p+�ͽ};��<fN�}�0z�Q�����AK�&���!��R����e�'"1�ʀx
wE��+
��!���j�66�S���慨���i#�t���ų[�UB0���@�:VA5,fq�~v�i��^�y�b8^�*F;sb�i'���hF,J����B����>m -͞�Ue�|�������^��K�W���8��)=�k@B��'*��)����K[A�[��2���������������Zw��G�lW0JӤ�#4ޱ���0�%1��l�GbYԒ���v�ޏR3ݭ�Fu8�^6�W�P������ْ�9$���#)�͘Mq�\m�Y�F-ܟ��voaK�Um��)qms��?�[^����+���+B>�oS��%\��]v2DM�c?�M5e��9N�
29���W��#jнx\��n-SZ��E%[����0�-&7-��w�/[�w�Im�y[��G�	�h������Jڄ�`�u�r�>���~���/�.��$�m7�ʂ��M�.>����VI�*-@ڽh~/�="���(�a��A�z@��ҷ��l��x��
{�D^�Q,�����V���f�n])VL�|��@09���8����?�q"Pn����n8�c��1If��n��?�p�O���M���fs�#-C�����+]Tϗ��:�Z[Z�����W�C"U�(��g��J�j��)ħ;�������-v����#,Ns�
�����U�����l�'���{N�:%�0�1��_=�g���B̦?�'�]�,�K����c��$���,��e�b~+Z��W)'����wu0�Al3�Ewp}��\�K���u4j�X�2�H�o����/$��o�RƀbU���t ����O�W��״QK��'O:�AK+��\���A�����%�y1�}��`.�2�$����֮�w&Y��G�R���nI��.�a\@�<�DA��m��?��P.y~��j�N��,�z��ZI�!)���b�1��؉����YZ�Y�`��x�
̡ɶ(��(V�r�BU�����١o��u`pI��ɕǷ�'VW��縻0� O�'Is�1����?�o ���@^��G�0F,?ZI(iM����M����Xse��'W{��m�=�.�,o/�o]v�� ��2�pk�R��d>:]H��l]����h)��+\XIƊ;`��e�nz|_j��{G_dN���e��
R�ܻu���'ud~�$%��+ *KB��6ak${wWq�e��jӢb����]�󶡧�g������Ƽ�Ҹ;��� ����k�]���%�c;�����8���I��eyY���+��P�HEӍ+��?�����CY��Dl)��1m�4����T�A��%�A��$1��js~��>��mG���{ٯ��(9�,���DJ�Y܀��%ٕn0�� ?��?��3P����0�����s,N]�:�/W�"N� ����ȳQvQ�{� ��3`c��!kjT��s���=�ɹ��gZ7Bf���,���L*�t�#6V�ve��s�A)�a|�ڳ�`��[��!;^�����E:+�K���X��Sq�p��.'��p��vj�]�{-�{l��,{cH��$a�b��v9 <QU��ج�M��7q��{7�N�E�{&�kܽ��6_��`2�jSBI��R5X搏x�V$K�Ч�/T���KM�5�P�����l�/��~n�#H��/V�D5]�r��4��M��:ٟ`��
c�NI(H�2&]�+�`D̉l���6"Q2�z����f1ځ����f��>�p\�#�Z�Ž�"����3��g�Pg���w|�����lE=�[vY�55��Z��d@�o6�u=��$Dϳ��E���ڈ��Z0�.��ߊ'�a0�Z!� '<ٔ҃oU��=�S���HE6\�TW�)y0�S��LG�P������<�T6S�^��Ѯ���ܿ���G��f�6�d{ѡ>;�KN+S��_�z1\�Ll��ܹ\B	��*ل��Ӻ�wJK�7>�TA;{�:[;�bp����7 ���<�*S��(�oV�"/�M�9��E��t;6�P�;+Lv���ȫ����g�+�y��
��6�����2^E�0*�샙Da�,��]Y�rҧt:(W>�&}ԯ��~n��H�Z����*�j J��=��ͺT��=��1�4��a�x~Ln��|q���x�߈�,��f]p@�sM��_Y�K���r|r8,��\�mw���F�.p˔b�_��uײː)�2S0��� �.���?� �a��aƗ�A��l�<"�C�d]��=�A��&�w�\6��3qF	N�3	
e�i*����6�G�l�n��˱�':�u��E�7H�jK3ԋ���/�����2�����	��ϸ7 �_V0��gn���]�m�6!J��L,NtWD�4��K�H�e�%,S�N1`����n�i����x�*E������ ���n1!����Wb�����u�~�=J!C?�hq*��Ç����AnC�f-�M<[�.�;V`250)�+8T�>�;������I� � q����c�C]�jc#��oo%�x�q����-[�,�戯$7�[w����p��6�o��$��'I���	�v�c���]6=��ٲ	�e���d��p���o o���'qv�ђ��m��>:[h�ϭ��̌��rQ�r�ge�G������9������u�\�B[�6���[��0��V�6��M���;I{�[�	G�c����&+�E�*5�s���=�
�5�~�\�c��a�W�Č�jVf@D��.�g UN?����vL#a�(��Ce�r1ovw�[_4�f��\������i���G��u8bk�C/��Q_5yS�jJ5o�9�%G�����h��-��~�=���:�ڇ��z
���M//Zr��;&ǒ���.BK�=�3\���:�=�6 ܺ?�'*ܙ�W�B�E�g�ة�O'x� D#�aZJSھ��7��5	30�#�穼T�ȶ5~��K0:��V6��ғ_ŃF� �ӇQ�ۇ����uc���UT}_Gt@l[��F���O�?�բ^@�Kh_|�tH��j��XZ�A���"J�?[�-�R���N�B�3�2"�{Rf����}�g�$��~��[�|>�::�oD᫈�2�Vw�q[{��_:�:��>eQ��.�YE�2�(�)�������$����:*�ާ#��V��3F��p̗<�	��`��%�w���8�&8����#������1֡R�ޭ���E������fYz|h���>1XlxVHYEB    cb82    12b0$;�.�F��pgf?'%N#��InV�7�N�0�K_6�4/AU�"�D�f�rw�Yq���R���u�Tf����df}J`�̲��+:��
��l�Ձ
J&����p�լ��ԙk[�:���"0�A��>�~0��~"u���Jld��}�(�!u�ێ����;�1�������.��.�[�b��L*oZ��͇U2�>��Oă�f���p��̂-�*��k������#R�wߢ��)����cj�sx����e��
N�^����eXC�u�+m\�s��2�;1��2�c��Nܯ�yg���0�Z�$�y�&��g^����rZ���Vh�j��ĥ���"Bl�&:o���5�W~�w��}����MA!��J�� `����(N��o2��:iKj|�g�xO�^>^����4o���u.�e7��b�۶���[��Jǘ4O�8�����%�ˠEB�310�e'���Jc?�^2IJ1�DEn��4�)d� �q,�`��\7C�֠�7�}o_ys�8Z]9$���̛rX��(	g���vLs|�Bɟ�^��4�#��`���Ss�l���m�$UZ�q�o)���R�λ�j��CPS�ٯ�ĳ��۬���`�/�����Z��;c��Ivzϛ�#�e"�&7�l�!"9��!�`�_�������miR�Կ�V4u��/��r��ѐ���b"���^\�㥥���������Y��`��FM�u9�ɡ�����W:؂d��lY��^ցE�m�Z;
��/v�\G����%L�(�W��$K�|J���x$�q�xI�>�I�z�Q"��8�����t�����1L�ά�܊��j��6C{f4^�S%�Y$e���n�o�c �9[����x����C#)����C��w>yPK,}��'���n��ͤnrV��?�� m��c���7^��k���{��DW�x��G2�C�څD�w��cm�V�_,�g��f[�U�Sw2��t[/z���֏kBc0b������}�r��U�e6���@=�pI;f]��L�z^���1	A��Ke��q��q]�ҩm�P#WJG�м.	0�X�G�]:|���z���`����gn���"��y�P�%B�j��6�^E�)|�(�4p4��x�؂�c�S���9w�����F�*�x�i^4�>^K��������sQ.o����i\��(Top��pk�81"�爗:�6�-����qP2������D�?U����-� ��$��ܨFk���c!!5�k`Qwi��L��,	p�[�*n����51$��D��¹�Ć����n���[ڪ-�8�-�@'����2#�] �i��dO]�e���Z���밓:ZUt)	P+E�l�GQC��8�0��Tn��AU,��]%.mܛ��~ƀ��K���w�ـ�xD<7�طu-i/��̲���j5����`���X���Z� `S�������y��{'m����0���ڔ?�JӐ(~|��*���0�
�L�PpHߙ������,��
(f���g�S_ݐ��3I�y��L"���� Evh������6� I]	%�1՚S�iG�)����s�W��Yd�A؜2~o�"(���֏���������Zl=���� �9ٓ辞����4�֠�9�ˌd�K�4j���D]3�U�;/�I�IT�\���lZ�`gY�]u�W�lS_�b�ƛ�����෨��o�2�М3�9>�V�ǝ�Px'��TJ����*+�� �R�2���p��Z�3�ϚD�u'UQ,�kk=��p	^��d��Ũ�&��oHE��!T���<�� �U?�&�8X��:�Ɏ	���ڕ)�新��u�A?͞+��eك'�L����V�P?�d9�ȕ�����_l`�bɭ�S�Q���,�GR���%�A�޾(uwW��pb����3j�7���j绍��K�>���	ܢ_���Ý��،7�ȑ[-�fj�,�Q�w�6�Y1"����<Ę���.DN8���^�@e��nT�8�L�-�Q���Ę7�x��|?(��0go�y��"N#x.SO����TޡÞ�rQ�cG��Nw�������E.U�D���;<b|N}�AR��W��R��Xb�y6���=2=�f!�4�4���^�_�8���'�l	ך�mdo[������z�)�����8�lwB�,�%}QQ�q���	Ko�,�d9�fR�w���X��+�Q��Z3P'�H��j��,����9�EGGl��#�=Nj���Y-�%[^r���&��V�82̠�#� ��@�  ۍ�'�,@�������!R�m���ѱ]�B,��ܦ���}t������E�S虛.	l=ƌ�>YP�9����Jhdcs۝�V��#q1�=i����<KB�+��	��?x����k8�W�&@� f���-�@S�W����w5sS�O�&�T�������W�-Pw���]Wg�S7w�B뺳��Ԓ�7�S�H�n�@�Oz�����A����>��|k����]���~�I���BI"XY�]��N��T���k? ~��YW؆����lK�@����2�Xzjj����`�R;�ֶw�}k>�>���K�#�2N�j	����3?���<�2
�KzN9nA�&w
���~<9�� R��;"n��I;�[�)�d������{v�#��N����B�8	�B�ZF�.H���V�~�O��$�W��hJ�VS¶|k�4zƃ��WE��Hk�jj�uTLzg�\�=��/��A�F?"EizR2w�̧{}�L��6��0L�WnC�^���I�06Sd� =�D��'�aS�3�����xֽh��K)�ٹ���y|�tu����� �9�k��u�׆���T24'a�l��/Ffb�ge^�i��u3gR��э�?�`��Z�ԡU8m��T4��x�y����ʲ��6��I�	�@�����s�*V���ϖ����c����t����F�q8����R7m�-���(о[xZ/����V���A��eȻ�P�;OM�{%5�Բ��J0&0r��!u� ��[��jL��7q���J5O�:���$?����=C���[x���d�^	��*)�	n��&�f�J{��*��-��e�t,^s���W������P�@�n���_���ʺ/O���-�p����Y��Ɗ��_��:�o��
 Ir�Z R��ҽ̎X�$���)�X��5B��ܷ�A~�H���!�M3��02� ��.�/�X=���B!5��A=�;ڳ��;A��/�xW�F�V@My�	�F�܀`X��ǰ|�V�4G�rQ�ɑR��
�pF2���6Ois'5��E�i�Ʋ����	��s��$��T7#�
2i�-���n��W���c��omf������o��N�E�.
$��ִ�*$����$��>uV��5D�h�	��תv6Z6�����MD��!qi��ar���L�3�_5�3x�	�`XBev����_Q9��S[f��[~'O��cY+Ri�Iz���b݊�9��Bh�G���
�	D���&��� �r^�I8��UG
���� ��3xeЗyF�����nW1�0��=n�x}\��Z󘚦<�/?���\u�;�Cv�hD�p�f��M 򉶾��X�»�Z�A煬L�\��TА�G7�
{E��c�lS̓�j�$ֿ����]P,��)5���;گd�F�@��I��pfh���'��b�:��@��Rv'o�lf�}�)?)n����I�_�;��p�����rt�����%;0���!n�)RD�-�5�F�Y��� H���C��_�Ѳ��D��4_L
y�|���ęD�f�~L�?2�E�*�qШHb;�?���K��T�$AC}�^\�^����T��n��k��r3�sNFu)�+� k{�9��dʎS�`Z��f�1#�NsK�7Ay�k`Ъ���!=�X8��sDi�U��[���p[=��d��/��qnP@FN���%��}����P�' 3��r\ϣ���%���"y�L96̻k��`��#�����zI:�%�DӋy��/���@P�����(�g?�m�ĉ%���}gf|� g��8�ġu1�.�qZ�e��,���fj��'y=%��o� r/�%�M� vu�6�æ�{�:�?2�T8�w��Y�	�y_i H�آ��Ѝ;Ś&ɇ-�����$wF��$U��������sVb(.������sz�h�qĬ�bcK)��S�p�]�|gǃ���d�8�y�q���z�<6.8SOa6VitOdڈ)�������j��>1���I:8>u:v����g�s������Z?<��޾'�ٜ�H5X�bh����>�������X��1����Z�$�����O���z��Ja�Nͤ5����R%cJ�G����S���U
�tuA��W�b���h�@�/�b��m��Q���@�((N���+�	k4az���M���z�m�kE-ȳ�e8Pnh��H�ݨr}�]XZr�9z�u��x`�����S�{T�����^gq��N�Ĥ&b�f_���YUyL͆��B�"D�TY}��0F�!��ч;"���ehf\V��x��U���.��e2�'�����)2vZA�,�di`����J���w�}������DyW����.d�`����|,m�Ԯ$��P9�<gi�aá9ê�'$\��U/�2ՙ�4�������mT�/w�
Ď