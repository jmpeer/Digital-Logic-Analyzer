XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���e��u|��$(��6lO��U1�7����c�挽���u���6�ׅk��?4�#`'����Kx��x	����TFxz��M��\Z'���{\�i�����5!��}N���,b�L����JJmW����:��;��0��C�?�R�p�Jlu�3��!Q�#��N�Os@uPO��UF��z[g�}�S.peҡ1Ajoh������D�m9f:�N�	��������^;�ED����w�Z�L��;�2�Y��;���O9+'{$��n`�6Tn�X�P4�Zv��<L�v��0�K���^i�k��8�
Xa�yx߻Nt�䞝�%>p�"��E����ԫ������X�qpMP���������g��[�?��A�oZ� ̪����4����r>�ܗ}3bA%�{"_�/��Σ�Ӕ��'���o��)�f�Fw!R��XU2�m{K
c���i�Z_r1E���Jy�LÍ��KC�b�8��V�g'h%QG.���'�?QV-ͨ&@�!;��Qc���+�k�ݥ�W%�j����]� &(����4l���ϑ��.��w���!F���Y��{9���m�(duv��U���h�iö]R�M�~.����D ����҉�vY>_��K�w⛲c��|��\��1�iߑJ��cg�����vy\e&(�~<���Ks:��xW�����i�q��Whٶ8�1Pya���$�~"�n�$Y��z
hXlxVHYEB    fa00    2950�&�xH�f���'!�&�bW 7��ʰy״xs	%q߮�դ$@�s�5�gF�sN���|��?*Wc8�mѯſsQ��9�4�D�N3�S��FN�py���Rn7v��P� ����.���L�߬��#��`λ�b�u����7�gjWyC�=���4?�p�oIA����CAA�[˯�~�L{qS�[CՋ(�w3�b�t�֭G���pTط�y4E��k������[��
�gBL�H^�سD��J��s�Q��^׶� �1���ED�ޫ*�Z}8�<�n�[��8׽�ፙ�*(�q�H�m��!�?ʒ��xA�_���9ݞD�#�A�y�o�_�kԏ���`O���}��0���������jZ�s��k��d�Ii:"p��{�刓�ؙP7������[9��@��T����Gzbxj1�h�ܨH��>@^{G�t�ޱ�Z4�r�׿���Q�\��=rAN�g�L��+9�_B�(�����5��T�b3��O��Q����-���dJ�/zL�T�
�0D����~_�Q�����m.!�L�wrT�!����]���_<:!�Oa�S (&��bO�/���f��b�`�8a��%sc�Ɓu��-������Ȥ�$�R'����a��*�Q� ���a��bB��UNH_#oᵶ f� M����X��	?3c��4���C4j�,0_�؝�$�w9#�HEC4Y�-��D:�y,��2�[m��tݦUz�P�r�~/\�[Pj�8�a
B�EC�/���� 6702�Զ<���uE�^+��:n�-�b ���N��et��j���x��x�X�sb� Ȇ�&o���`2����半5�c�9p?�m��:�i���&�F���i�%	ڐ�A:Dh��n�^s�Ӗ�VA�Q�,����Z[�$�����B�=�L]�'���i@�0k� ����	G����y��D����+�c�+�b��b���G����|��X7�9z9�y�l#c�({o�����j�"�ȗ �UdYP2�DS�C�cTGt%Bc4ˇF���T�>O��� �?�1�}��؇�i5ڱ��/V�La6H+E�i����?tՂ��O���9J��g�Vk#?����9M�S3�F���vU�=#Dq�fG����oV�c��iǶ���I8�����!�s���&,*y��fW��P�X�6�0�c�]���]Z�Zm�w�>jx��>���b��&�wUp�<'K��`�&̏�Dw��l��eT�S�/娡;��Aı�6ET=cF�NL�����A��BqY��M��udũS1Yx�`-������YXx�$����I�9�������t+���p���
��1S)���wگD6-@���/�@���a��'����L��R�:@.�%�>�Jd�7����(�$�Ǘ>���+�<l�li8�g�T���/\�|ߓ�C������|����mY��Q�;��H&qZ�r� Fkb�:��C�����jYp�QQU�F"wT<��nMo5��6�8��"�<ڝ�^_+��%ueSC|���9#���XYҴ?ǡ9b~���F_�f5�:���m�u�5.�%��Ԩ	�9�<.�:�[-�K��_��2��)�^>�sR��;K�%��q�����Ґ��D]��-�����0�/P�A��d���xk�1�w�i=b���l��vWt%i����6/,kGuo�W���ޖ�bW�1%��;�\b��=E� �G.�HP`G���U�&cU%\Nu��Z٩�g� ��`=W���ՇN����
�W���Arݦ_'����\��Ũ��+o���
��Sh�@x�oRL���o��̇^��V��6����?*ڸ]`T`�,%�a]x���q��)^Ԧ������?�9�e�a�,��+����� J�.I!O��^��4��j�ǘ�����=N���^�[M�I�e��֯~AMO���x�],f���2���ؓyYmu�tN��W��ٝ��_�C2�T��:=3�fI��������:�E��	�2ݬĈ�{�̉[�T JE��6�r���{�n4�<
Ih�.s�kN��Vr�����ܣ�W�)�ǟ�B��c-�g�jK�ĺ)�:�e?Z�A$�N�2ۨר� $�h��G�d;l���t���x���R'���=s1+wxE�tk�h�����=�z[�O�٤�{_17�w	0Л��3@��+_����%5���֖n�R2����ڈ�_���8��Ad��3��	J���I�"����Z��/47�@BҺmh�,~L�8�\�7Gd˿�+��m>��}x(u��E����,�wc���]Hr��E!6[����Z����b�44����-F&Ef�U�a�18��՛�k�>�Q?`���ϼ��U2�Fo�P':�E�ӌ�?�.�W��C#_�dRh�I>�T1 8��"\��Q��E� ���~���<!+�P9���j|d)��V����Vp��
5�		4'� X;`mv5������~qL����m���~�cyw����W0�*:��vr��؀6PO��C��̘H !�P	M������r�B���Q��-��$��0Y�j�8Lih��T�=M�'��Ny�/�m�d��Ge-��ܤ��Y�n�i� n<��y˚��K�R2:��;V�)��t3}�X#s;|� �h؅rK��o�W�ۂ�ӟ�=��8�S���K �1,��NCr��&�e|�k@p�:��x�މ(au5�_�a��O0'sӂRߤ5��,o�GM�����,ls��dɇH2����Y��#&S�Χi��y�9�����1t�d�E��@�@�y��ц"��A�e�g�y�7wU��˂��6j�Zp�� �.��>w�$�!7���*�j;��]*^�Z�pE��9NsL�+.�c4@��8��z�ͷ*�
�5Ix��C`��W�^M�I��ZU��gFnb�-V5-��d�������4U�����?��Ub^ۜ�P�=/%�@��`K�����FD�M,<R�[H����x�|�P���k�9۔��?�^ٙP�\[�rE��T��6yj�����~\������,�GW���df�Yl�*k��sg,3]���q�;�}'@��d�F�7W���
bY�t������� Cb���>o�,%�.�V6q����7�{s���Ev!���a�Bi�֏�63:zX Y�\<�P��c`��[U��j� �q��xd��gD2��X~��r��0�Ȝ�m����H�P�w�?���9^t�C� ���"�0jA��L�X0�������Q� 
H��4��[��w/y�V=����Y2���>�g�O4�$x����`zb�ͅ٬J��
��_�H� >�k��|XGB��Pk}$)6B���P�0-��A8�7H2��
-2̈́+ |^�;��T�^q��c �졾�w	$����)�A�����X�"e��N4�b��`vfy�2�nl#ž�G6.:��'l��p������*����ަ���l�XJ&3w+4?SQt����x�����೾�C�H_
����XA%~���s�FB���}e�A���a��|��fez�m	?A��UKk��z.g����b@�&���)l�뿁��ˠ=]�/:+�nӘM�Cd= ��F�t1"�?ه)*��鬆�P����E�5�Q���2���#x׈^3t./�N+`7��6������)�{�vط�J�����T����p�(��2�r��
���1����휭l�j�I�Q��\���M{��Ꞇz1T�۫��`���
�P��=Ϯ7��`pO�j����)!���z�b�\oA|w�2髟[��>��h2Z����؝F7���I_�)(W*W�>u���IodT��{����r6ų �����!r�dmt{gʭfm�Y�����&�J*=~�}�W��m9?��\bݰ��S=�C�;k3V
��}���6���	�Fm����v?r�PKAjs� "�IF,q4�Uz���,b�[r!��K�t$�_q�ʴ�B��i�~.`9�?����eM�'j�;�Y�I^$�8[���eֆ�;�5t����?��t�w�p6:é�#�F���3	��,���58h�$V����<*�SW��]"q/Z.�q���3�ƁR�~*߇��}M�e��O|�n .�	��&�k�]�u��\{4Z>�(��N@��{� �x�9h�,��Y
�"O־Oo��m�ϖ|�h���n�/sxf�5<Ļ����~;�n���~�����Kx���F\����7�޵��7t�1#��~r�S��<�Q�7P��q�^
�l>�����t��OCj<�ʹ�Ab٤v�.���Xxn�VkB�����xb��Ƶ�X(���@"u�s6NC	_�\3�F����*eM��9�<��X��#xE�\�V#��7�%�"h>D9%�	�G����̸``�*�M�U�b7�m:�Ч��@���S���*_֊A�i�-�F�ӽz�� l���qb[hp��u�� � qI�޹}a�ɷu�|@
����:���ɐn���g����X_jZ�g��G>o��d^���ͤ���&4�����7�K�4�1�!�m���X��!��[���������5r�������=y�xya~D��Q#[i8��.��W��O�bd\1�x��O%�,^��|X�Xf������s��Ib@i�+��B�����+r���7r��������",��
�	Sh�@�GÇ�U��ءs}����*��m�7t���Q�凒sR��)��;X����6߯� 0�;������<���Ŋ��A�:/���M�

��f3K	�TY�K�_	�����ƋY��T��k{���.�QؔDwi�4ۖ�>�����T3�J+�Lz ֨�=^58��<��0[��TK�G����
���i��~6�"�_��O�Ѱ� qI�F�g�Ӌ�q��S���(5�/�B��L���C.+e���C롢.�c���`��� m�q��ek7l
θ�o�wm���Y+w��g�*e�cT�l��$/�L�H�����zg�Y���6��r�&JJ2��ű�:蝂{�gB�PP�۶���]-���o����b�� y����b30�Ӿ�t�@�k%O�k�e-�3�a¼��(]��|)��x&-����!O�������I[8�ޭvݍ�\f��Ñ���*����9����Wn[��ο���4��B�U�e,1�6-��%�r~�(y ���'6Ì��U�8�{A�5� �#r�q>��;k��:���7:������H��h;NV���v�1va��Ȱɏ�6Ŧ�ʶ�؇h����XƱ����OLZ֎����f�Li�֫i���v̮� /E:�C�s�X�q��b�b��1�����TU
˔s�n�`/�(Z��!%5446�WfgXՆ�GYu��1��Uݍ���>2=�v���?����O��[ܵ���m�;1�54�g�5p���Dӊ9vx�}fW�(� ��x1�W*��0&y����+��
��M��!�Q�N�c�<����1�A�r.$��+�+*�+�>;�&������2�L��5��Q	����Q�ſ5Aax��0R��Y�4.���F=�/'��(aƥA�j�G�39�fƀ���0C*%�S�m��OU�Z�9b/���5��*s�^Q�a�+o����KR��2������oa�V��<���~?^�W��jv\2!!�S��5�96�E�F��A<���?��w/��&���2�p�[�e���ւ�7ݷvC��9T���1���(`,��Q�#���q~\�f���&b0�ro2U�b�M�?S����]�|��*��]�m��=� ���ъ-��|2&>�^vx�+iwY�΁�:N�l��o����@yH/���"��N���D�2S�H����OX�X3�x�&�Lx�2s�`vw�
�!�;n���M*�Cg�o�gP�t�}V��Nv��O�,1[�_Xh�(s��;R'�<�1���4ޟL}�<�m�l�،#�9�])�8�}m����
��&�+���垙�P�R���+Te�j��g:�bP�nS��(&��u�W�Wbd��4sa�38K���߻CL]_�!�}__)�d�M��rnߚ*��(�U������Q/���ة���3g^m����v�G��^;/��H�ͨ��2u
�y�G������ΰv�6�"�шtJ�G��V�	+�5]܏�+̩&caU�yK$���LM�d�$e�i�.����=��<��������wK�L��r���79c�2� %�\0ۛfY~kl1�RSCۿF�w�V���(�G�#�\V<��;��d�z�MNj��򐳗慗E�qC����j2jk%��<�8��Wg�`�KZ�rZ���0Dv����|#�-�v��ʸ�r�Fr`&��(�t�j��ݾN�u�I�U�d�ƽ���=�'9��׶��j	ˬV�M�����s�⩱��)S`m�1�Nn�bӖ'Ҋ���
d99V0�ݸX��/�UKBKcK�����\�a"�!W�cR�f������A�����-��!�k�
�����ysV�4GlK
�zI��n%���C�	P.�.���+�&�[Gć���[���o�B���;.T5�u�5����棎�R]���!(ѷӺ/ܫ�ρ*`\a�@�]@�����"��E��NSZ��:����t��oG�3�,7$�I큦�:3�@��w��z�2?��7�i?	>_�y�Q�^ϕ6�N]0w`?�ݞV�9����f���~�ox�s�#�%m_�I͖{�KĪ���!�yz�?Ǐ�u]&�!��ֺ��u�ĺz�
�T�mNP��J���]ǬW��"í;��?��Z5�n5��*&Kw��W\��*������n�M{��VMD ������aPal2c�{S����/m3����D��C$��h4NU�t���%X��v#��U������x�M��Ç��K(̳�a(����F�3�Z��xRVJn{�����������6�Ģ�%n��m���I�l��2rH�����C!���w�v���{�@1��=	Te�/fTt�5�I�vU������,��Sa��>��j�^ �H8��KbUq-t�er���H�JMHt�*ƹ���=�"�G0g6Ŗ���$���G=+�x~�ﶛ?��왋J�M�AR�g.�HRɨ�*QKE��2���M$��h�F���̷�<��ᗪ��(�#R�P!��BY^?
��BJ�<�}[��I2�#��hO���2>���9Mb=��\܂ɭM�E��138�E�Z:+n���x���$(�0Kq�ׇ_�&�+�R�v�j߅t3d�צ��&"o^3����F���qG.�q���@�B����p��tF��<��K���������e��|������c������_wr��G�P΢QH���	��t>�B[�ZZDA����H�4��C���B���|p�y��
�v_Enf���Ulp����c��$L;��PT�q�ϸ�r&�@q.�g��̵h�9�Y3ϣ�I��9�UO@�U��#���1���pQ��~f���R/s۩���d�A���p�T�]�-S��ՁGy�U��kH/�u��Q~�9�`����c��l�h�S��ý�Mzz)��4n�^0�� Z*���k��A�r'�Y9��r��:\�ĂT�h3�`SIs�9��i1�\�U�E޴a��WN�d��4q6�tEg�t|�o��6�K�����@XX�0��V��z�����mms=W*'n�u#�*`�`xR�Y�!Ed���DYX�f��ձ��}��(4����[_����GY�������s��Js����h�?hyΈ����f��S)C"���	K{'_K���x�������ox�0�\yP1��j�g����y	_d��%A�Ջ��jT��i �CK>������Ʊ���`E&�A�p��8��4�(+G��Ci�a���ι�P=�C��2w�aGn~����}��8A|ڎ@m��fK����=���;�3���o�fb���*i�u{ǃg�)�A~m8����>g�O����;��F�.)��ǈo^_OxϞm|%���c-�"Pن��3�L��j���ץ�2Q�� ��D�����?7��)��}�(����+�^�):ޑ�׵�=��Q��R��H����:�)y�!� X%5%��g�d��,Ꞟ��+,�"2�S���y�-�'s��5���V��NK'8 ��?i�Vv�\5�E|A�&z�R�	���#u<���6�ɪ�_�M�Iݎ�J��6��{^�KN�oo�����T���ot�����ƚ�,*��z��p��	�6U^����:��U]����]R���,%N�^������Q���D�O� ��o��W�,�l���MN���/O���$�Y�NҶv�g:� �]�L��u/�����nr�\�A�%fDy|�����R�K:�-�Q�X�������͒7��3[VipR=�o��(��%���Sd��=��;b0m��&�������3#<&����G�S8�$׬�B���/�4�BeȽ1xɥ�E;G��e�y؂��"����rK��y�ƚ� o,��y�a$�k>8s�i�3�{7P���K�7��d�U r2';&�Am���8^ M �k���#���@>�=��zq�ՆybtӨ�)����k�j�f�ݐ\�d� ��|�����*M,�֢���lh16��dLO���@"��eHz��
utA��Fl�/���J�v���*��uѳy��T�����ز���Ϻx����$��F�|� �橎)G=�+ꓐ�ː�c4O��S�j�@ژ8!�|U:}�������e�����몠��hMY�+k8U�{<��j�Z��3LR���ӫK3<Fڡ}�S���N�Mp�BS�Q���;3�l.���&cGO�"o���`W�2���ѐ���Ő��G#1"F���>"���	����}�5�K�I�i�&Z���dt�v��6�(͐�'��$d��H�(a�C=]�SX+�Y �fa�dD�]��ǐ�c���e�N��8��&V��=��GCR̉@��V���"_[ 0!O1YAfy��a��B����K&����0�»�,�=+�qu:�jl�Ei�A�=�!Ad�R��R�[�\B�\�����2���?L��%*��YT�dQŬ��N<�e<w����*��Poc����t�ٔD�7�([�5+%��N�P�S��z4�e��� �duN�U�`wu����]�3��9��6
ж��̱���f?Uu���������v�p�L�V��|ƪ��6��!Jm�;!���c��������v�Y{p̣�J�o�K��D��k@S}rbۥŞ�XEl��2H�ˌm��ք�]EVq�����ΘXh�Tp��'�E�k��ŕǖ2��~a�}�Cq��v��	֯�"��$�HO�=�x��A�K�z�.;ڶ)�x���ť���&,�p*�K:�`��n���	���[@�TS��OP��]K�� �Ugy��C�yg�$��#BDL�cB����ԉ��[����}�J�ali�;ܭ ̀u��.�����W����V�e�,��asQqc%}/�_/w��v�K�dn�@f�T?�Ѝ�x�&N��8�~a�^MIĖ�Ve���Pƴ�N�E��u����mH�����n�T�1h���K��b��������E|u��N4"n�����)���Ӳ�<��r�WaO!��:s�1��w&^�hx������+\X�����1��5P��LƖ�:\�d��L��� ]��Vh	+PewJ��v'D�b��4UvDfv Am��i����H>��j��E�ʌ�aP&;6�Y���"�	��4���+�-L¼��#�#�^욏d��$}i��,�}��p��pS"P��^w(J�Yw������r��uA�Pts1}����yfz�$�謙�[�d�!!E����R�N�ذ��١%��*2�a>IQ8f��`�	�!Ց��ڽ�x���8��n�իM�a\�kڱ�_�iG~�2?إ�BU8}�o���
"���K���9k�o ?n�!ۆ��b����촩dP���o꜌����c���E�PȬ7��x7�vm��>d(�It�Ӵjx�|�YMp�"-�`���;�����;�IX'��+,k�垍E��=z�1����Y`�K�\TD[['#n�
Sc��m�̷ݛAwG�+�{��D�QR��K*ptL%H(�4*�u�8�B�`�m�9l
mV~��l��V����'Y�cd�e��E�<XlxVHYEB    fa00    1e30ܤ�ʧ�
���B{��Z��"k:���9y������?�Q/���e��`�j�rכWE��Ǳ$�R���k&?��Hb��0�E��>0�g)�������6�UG�B�N*ڸ�.��^Us�̈Ci�4ƌڨ�ޯ`s[! 4�G|@���Qz�	�>��mL�^ߛU��a|��=H��\�7@_��{���9��ܷD��w"~>���m��"����RIH�*��Z�V@���-�P�-������ .b��e�*ar�;��'^E;���Y�+
U��.t���������]��Y��tK�+R^Fu!h`mjs��_*�uzs$�Z�Y�N.!�E^�x .^6�C�^e!��Q���'z���!l���yC�i�ry���5�'2��S)BM����x���gtKΪ���T��C�SJ�@*3�x5q>,��`���>��3ۋ]W	���D���{~�q��,mVQ��bM|nGɅv���
�FpA�$�J�&�&.�U�ò�+�Š"P��+`��&zi{�y]̖���lه����
,=�����oh�k����Yzś�&K�N�����[��W�e=��g�|�Cj]�>�I��%��-����Z,^��ź
�H�
\�@,�x�薱��s����s��J�WI[m$�Q�+Å�ɃH]���^@�O<�!o+"O�倲eJ���/��x��ܪ�C�<�AS1D�����M�,���������sV57����[Q�`	=A�2���Ȥ�/IW*��� �y�E)2���E)(QU����g{ۤ�G��p(��ʸ��$�b�D��5�ڛ5��=!�Xɥ���Kf���f�i��t{���(�S�9�iFf��:�����р��Y�eD��Z����cQ��D5�Ѽ�m��
 �q�e�#� qvEt�,&�,ux���;�l*����ԫ3B~�H�-��C����5�㰅�h3x�J�u�J;�����]	BV�c̶<��F�ZT���K@w��d���==@!��?C4Q� FF�m����V�V��0)UO5���mB�@�{�29@��K��D̭�����9�n�����yJ���	_~^x��,�`nb�������H� s݅��Y�Wi̹����IoI~���W)�:F�����ĸ�R{}��79偈����g����^g�9�D�s���n7��_n:~���AwG�g|�uZL�כ�P*�mţ�\�
.?�Emj@��OU����{iM��g"!���n3�N�e��(:�!4�O���ITj%����Ȳt���s�+��k+uF3�$�R�gU��k�ǆ|�k ��5ħ�1�	����ay����\�{=:�
^��0oF��t�c�����X�>I���=����L����
������ۨ�I���ڕ1�mI��=x�U�܍{�T�o���g�Z��_��B�����Y�M�'4u����z�;�H�(5BC6(木�V �{�/}}�d���Qn�����,��N�+���%��[�{ v��'O2M��?x���B�亗m`�Z>�F����ą� !\0퉵��V1���t6��Z�сT[��;g=��`8|w�G�ϑ��~�v�����&ċ*VH�j]��ˉ�����my�'�3���+ i�s�µҶ��.Ҍ�A���X�D�y���]���&´%�9�O��N���s��zlHJ�όm/��#�-z$'6�^���[$�G	NF��쀩���S�?����{��u��8��Kn�kf�V��+,t6G���������iϙ	��j!4�n��SuNx���+�&�da�7'�(�f\�G����@т~4ݓ��iQ���ɧ���C�ۥ��R�_�����%,S���tG��LF�rU�V����dѝ��W�FB���Y!`�$%g�Oܣ	F���^�m!�Ɓ8�J�̗���^D�1����knW�@F�`1�4���H��W�*g�X�2nu�w~�������,��g�w�W�N����tN�/�����Yȿo<LYdw��5-��s��C_�۹x�i�	�S��}�xFVO��c*^�4��{���ї��+���R_Q�h/�_,=oG���'z�?���i7�����k���
���� 2h|i<��i���M�]i��q�3w$���% 	�������H<�Tc�s�Oփ��q�K$�.�	�eɏ�����/���$��~�UD��j�yFrJ���3�5������=4Q�j74s����xc�i�(@Z�E�E�@��T�h�I��8�I��5���f6�1{G�c�\�Q�RF�j�г�_C߿�X=V ���0Y#"E�\�:��\�!�L�L~��K�t�k��f`���I�g������N�R;=g@a��X���[��3���䄹�v&rؕS��s%M�^Z5����x�C�&R,Nj���}\�OՉ΂I;t�
xr]�NO;����]U:�๥"`f>�H]�jط_�m�ͯ �m���Ja�V4$�_���X'������GqQ�m�|V>�
�@7�����O�m@���l��y+H��.i��T��#�=D3I���
�n�M���wv9	Ft}�8怎���d퐄u@��FZ�����:����G{��J��恖��#L���0���x�RqLj�*r%·E�j�h^�b�>͒!a�LWN=��Lz��|��-�D�G_{�g>�GF��d���pOo�8�(Y�K/Jj&)����k�qukb.ޛF3t�jN���p�ɀH��9�����g��,�Aڿ��Պ������6;B ���B��KzުGB�&d�?5\ ��u��L7̽N�]�0T>�-:����	U�v��f�&�%-��o�B~��,�Z��]����7WJ ��|��z���;��K�*~��b�"M���EN��j��#���o=���1a�(D�րg1� N ̏{�Ǭ���k�N����".�G�"�� jN<E[���Z���fő�t:�T�Dx;gE���ζmN�[���-�x^�E�i��xMaĳ��>�zX O�ڪm�!�CJK��k01������Ƃ�t[�tBS�N/�p�F.T��u~��G6��`�|{��ud�#���U��%X������Kϥ��~ς�ۿ��e�:�D�8q���Bn/3.p��|�v����/DhF��W�{a�-G8�5� �`#+]��B��b�ZKU��Op��z�-�W���X���@��Q(O ��p/mvo��]8��\ꮾG�_N�jT6^���8 (T�U��	J�Wʄ���0sse!��X5���މ�mO�,�܊�؊o�4"�����<��P���ǋ�Ry9A�6�UG���_����n̨� ������B2�K��O��C#�I�� �y1����v�yǇ�Ua3�8�+C!�佻�B�Ļ���B�>H ��S�A0*��QXlF,�,~k���>�.a <bd�����f�{�͍,}�'����y��_�kҙ�d�Y��9����H[e�C�75����7{ϓ���!v[��R?!�3����QͅD_�i�8�./n�I�W�����p�\�.���*�M��������>�q��!�v#J?���ި'`-P|��eǃ���%���E[}H���K��n�O[�X�5�7�����(��$Gǳq�ue��]���z���>���d� �7���[u����[X1�7�h�C'�?�rDU����i��}@�w���1[`	��4�Ⱦ���1����Mi��=/g��߆A��y%�^���`tUʤU��F�G���` ������>E.��0Oo���33�m2-�J���P�G"�0e5�&��A�=c守v��e�My�\�4M�5hA�?�b�W��㺑 t�'�;:֒�!�O��sP|b-��h`0�+e���� ���h����[I9��I'�)Lgu��\a�S�=%�u���OP*����O >0�:G��κ~�qk���{�IR5"Ǖ�A0H0��z7�����\XcCQ��גٵ6s;��AH�6{�N�ӷ�{����U�5S�h|5����0��z������ �$"̌\�L�К��ۆz�g���Y�*��M��g���H?����x�5�ی�r؃�]�O	��UcAK���ࢼ	���`��;f�x9���cq�������"Pׅ���x��髦L�e�Q�U���7/�#
d!!���(^%H"��$��z�-�t�zk�\��ѵ9�y�R��G�ua�p��=?�ǂoP��2A�tƹ,6����-��0����_N:�5������+�QX�����DL@Y*U{�#��p�N�|�'۩��
���E7���7�C[o|~�Inh9���c�r����O���Z��O&�����*z� |�.��JWa��p�i�C�A��s�Jԩ&�R�$^/�r�U��t ��]�h�<��,x�ש��r�b-ݳ\iM�k�ߩ�Yf��x�\�1뻨ޝ�D�X)�C��6�+oaL�U�͖�
����.�r3c,���T�G��J��=�Q!22�⧞b�� 7�U'�W�� �:�^�؇��4��ٟKې�"v0XY�#`��*�������w,�8JM
�)�)��ۣzl����ڑ��K��y~���S�x�}�ݩ��٢6�	#烱E������@F�k	�!�ʟS�F�7�pB|�Gqo�kt��|)Չ�x�Ϥ�@΅۶cPi������;a�~n8��L���9}�@�/�+4�+��An;�����������V�&#�QgJ���i�R��-�\� �F�|�Չ���	�o��`JY)[�p�N�%%���F^��2�C�0A��6^2��[�Ϛ~��縉�]�<N=�P�`/�%`sYx��ÜD��G�4������71gb��� �K��y�[9lm��r��l�c�n~�����h��*g.�z������a��m!�n� L��g�f=p���9J�1�����������rc(9vo�H>|O���9&�����9��i�Y�iy֚LӾ�*�,!v�Z��E�D�9�4ت�+a���P����㴟n��U�+�7|x�Hwn2~�!�2 �a�F�RHg ��������|.'���5!s�Oz�.Ǖ����3QB����n@T�M��?�L	��ҥ�㻖V�����o�>O�d��.�ʫf6eLS}e�a�ב�>�Y��X�L��Tt��]���[v�?#��B��<D�^�$�LYt�G�r�d1�i'@����)"#�M��o���s���X���'��s-v�L7V<��<G>�E_���K>Y ��ږ� �*��Λ��r��ξ�/������ҨZ&3Y��ݖ��2�˖���"r�o+��|6 ��"�Sr��ŭ�:X�!~ڟ�� �*U=l+t��Y�A)�8B1ۣ^2��5ӘܧrDx:��?�X�@��Co�LP�澜��́;��//R�ja��x U�X	F�-�+�yل�6����m,�}M�cPwF�6�/����߉q<�T�d˜��>oB:�Z�t�a	��`+���,��4ܕ���Ќ�8�n��v�W����o���qjR{ٝ���P*Kdu�W3��l���϶����/��ސ��
/�����S�8ᑧĂH����B@��wakJ�.���:{�vN���t	�mnr~���!W�/=UmQqMz}�.�6 [�e�G�j��&�}���r#�}�u�����qo���S��:�cv?�Sދ��AX]�e��K(��/���~���/m��Ѝ.�E�dwbͪ@"̃��d��
_J#6�\�	���cu͸Q�<1)d� �W+��~�F��K������lz�ŭ����aN����|p*��(B|�A�`�I�L"�}އ�Y�l�����/Ǚ��g�4�\��h���J}S����W�����SD�ct�+M=Շ�=�9?8�dkmWk�3Yv����2⊣��<Y�W��Q-����ך!� ^����Ҹ���O88��D(�%�UK_E��#M���	R�G3	�Nd�z�x�@��O\kLd^�`� ��gb]�QK�h�֕E(~&��_��ױV/�le�lF以�.��]�5�:$�'|=��4��վ1��o�`!��$H���B8��}��e���|V{����6��,�_��P�
`����I���ct�\[{�A��;0�����
;~�TP����,X�Axx�7�
2�,|�u�1��At�_#�{M��%��?��N�(ܳ �[���≻�����Wɕ�u���3�Ƚ;ҫ� ��&B�;]�+��f�+���Y��F�������9"ӑ6~`"�_��W��E*�d�%G�^I�+0�Z�&y�C�ycM���_Z�]�������j�>�������y�
-3#<;�3�O8%��e��������l]a�s��R\�2^c�<��PT[���n�:K������ ;�=��6Xď��jZ׃'����������g���c���e�C�:����lJ�4��	Nӓ�O��τ��Zv+��Sm�}�·]�πe�0�˕����ܥ��{���\5}�4-��څ
y������U�<�Q��1M� *���X��}��
k�d+�����:�V�:>i׹�P��-����M��\)#>�5pz�b@�M�:�21wn|�qþ����o���^���P��DqJ�u@dr5���>��~��֩�?E�����&Ӵ(<�cP�V�����9n,��SBcNѻ�.���%��$,�Ҹ������2Ai�����FU���Twq���@�&ɓ>���+�}˴0z��n�|��6@��}���#Z_z{�G��ٹkW�JZQ
�Q��c�Lک�ݜpo�E2d�����&����, t��(b�N�u��I�Q�"�|��p��v�~-�d�p}gT� FO�]c�1q(�a�;�78�D��*�U�h
�u��P87����%�,7����}�R11��'p>\D��$��]�� �8��	{��R�eh�'��bՀ�g�ϼBC)�I�`�����5�o�|�ڮ��xq��*�ld&q�,���r$D�ĲnAp�Sj ����i�W��I(�}Yf�L$�&aqD"�����,u?ø8���6.l*d�����/��P x=�c7�-���!)ބ	��HJ�>�&�1
ؔ�W��,8�Y�g��ط����>��f�=�Z)Ai��$|��[G��;��-��J��\��Bۢ�,#��Ƣ_&��_��
zޜ&b��;�_'�dx$5��,; -ZMk����	��(��~�k���Q�F��>�q)h�G�W����z,S50�u�s#�S��d�P�HX��9��������Lh[�^�Zc=P[$�CnM�{FJ�׸�N}pj u#��;04mV��]exOCi��v�5R���5cyJ/�f����z�Z2lK�ޟ��*�^=����C�����S�σ�R�[S�Hpv3:��h�.W���q���v���Z����f;ܣ�u� ׻��	V�춨ϳ��.cE��(�w�����
�Uc�d?�B$�:o��k>5a�� F̴-]���7rŌj��L3lH�����7��Z��XlxVHYEB    fa00    1d20�_RS�pbWg����^�wմ�.Q���CTG��f
S���F�'�;����N�zT�n+�肜���}ߙ�9�]я?����m���ꏃht���p�"wF݌���ۮ�؜@�δ�����\����zM���Ui�	�²O.Ԥ�g�?�p���n<L�b���)"�G������	Oo�i����|��2П��®pW3�RF��Rp
��0oE���88���D�9R�1��%���t:�TY`�AD�΢� ��DrL�JdXì���g�Ci�5u�{�Mс%C+H�g��f�^+95�h`1��51e�\�u9]�������H�9�h�D1�;����A�+��W{q�rG�/���swX>�]�?K�m��\��v^W�-�C�Bݙm$yC�ο�0�d��`��"�ѽ�����VcJ߫
������4�=C�؋�7�M6��{y��}�o��H���(/?����e'"�9�}�/V|�4�y���D�թ�#����S��@��ҕY'�;�L`����H1۽b��{���s����3la��~����ά��Nt�]0�~+���e.}��P���;�Ҟ.����J�m�e��1zr�;�)��{����M"W��k��4NS���h�l8�:ܩ�^h]� �Z����I,=��8�{�id�"��k�:w�m���0,w�"�ɳ���z䑒���1ĸ��{ʍ*��ѡ�ޢlxpq���+V��a&�����ٷ^H���r���|<)��~��.мd���piI�d�G*ykz�u��F��3�����'��8jӼ۠:-=�>��'��|v��Ц�O�%���U(��GЧ!X8�&���'����yc�S�:��դ�`�S��E�;��iw�_�
�ƼQ<�mCqEai±pͱ�P	��)�'�UTqms2 y��#�#�������p����^��,�^�5;���8	��Bc(�o�"n�*�Tk9��QX�b ���p~�Qٳ2���0�:G��-���M)i&�>nϾ#{���N"F�A���.Y �?�nfmRg�H�c��|���e}k-'���U}��6��B�T��2gG�ނP�������蛪b����z��UB��0�H�7��'��7���ɧL^]cK	��z �=�?E�D)���[��ѯ~Jߚ-���&\+��:hj�ƻ����i}
p�d�"��]��E�1B�ɑ\����{�/��]�{�z�m����[�`�3+I���Kf�l�(�T��³C�k6�V�bަ�WX5�<U�*}�=FK�|X���_��Ҿ8�6P?�OǓ~�{�]����I�Maoղ��r/�	#M�����8ƁGr��T-�܊���8��Wh6�H���sy������Cǹ���>ҽ�n���N�����
}XU}�3g5�|썗N*ۛT=!L���_b��D`�:��!� Tu ,ٙ7��ck@���n����i[����s���V1FIb5�1O��g]τ�~f�Y�#09�������64*�uYX@]�xi^x�]ŵQ���V��:J��U��*�Ҝ��
O~�e��b�S�r<u�������J�=KK�@��9��R|I�ۄ~N�o�ХH/�����l�B!����a׉��{���}:�}���&w��¿���R���Z�/���:�,�fN���ڊ�\H�������	��|���2�0�7��� m���6�s�����O��塒�܃��Y�f>�/���gj�VI�t!T�y���O��s��)��=�)�p�^N<9Y�T�ϟ��o��PU���/\-�qϔ'�ڤ�
�o4[�z�m��U��c�y�SZk*�g��]LS�B���g�?�2�l�p�^�w
,һN��Ӆ� P/�V�oq-Қ�A��گ`�� "���?��ӫ:^0A�Ugor]:rF������m����a{"��/����� )ݓc��3~?]n2V��t�҈���9v��嶲��s������C�4x������ֺʄ�A�+���F'���^^����+�\ތ�~93������gB�S��q��N���W9v�N-[�^^r��+�5�u���&5P��8v�u�	 f�kO���W5}F�����(*�e��&	�u�+Ⴛ݊w�ؼFO���E��&�/C�oԗcb��'G(��b�@��VR�#gl����׮�3�Lz�5�a*�&^��F$���Ѥ>(�Cb}>���~%��9���h�|0��k�������*>#cx�E�XF	AA����#�Ђ>�!7Y�N��E�G�`:�;�9�-�pE�\��Hl6)^�+������<3����rlk�I#����қ��"�
eAN�#�:�K���X��	�3�]��� +9�>7���-T�h}�k���p������瓬�)����g�yўKʇ���P/�.���z1���� �QF!�@����[�Ă8(g�Ոy �XO��g>c�/�r'0�LM����&�`�Z��ؒ�;�wB�6�wXY>�0.:G��'��)l�
�}�,/7f�p9����ss��T/��zI��������rD.K���QX��+��HH|�]�jz��y�f"�/�E��O�����`�.�hrH�������%��k�B�~�Y��|�������[�n��G��b@��- dL����)u:%:���Ur��QPp��0�ؚ y�&>Q��H�K��A�F�2	xG��'ʪ\����zt%��`è�o�Z��L���Q���1�K>����ׂK7	�D��٢�+�IM��Pǉ��u���,|S��)y�r&�Ǌ17�=��P+��uve<��p�{�盉Ke�D���.&� �UHM�Q`����G�!�b�����-	-22`W���� ���(B��B.qᦙv�o}Y������ ������Xf"�Y�S`'��G5+���a��c�gH�p�fϰ�}� �Z�Wx���t��Z6_�-{-�X B�tlg	���fP���9Du��$|ޡ�-���g��Q��p��HW�M�v�`�ʆ%�\�'Qx�'��M�)`:����; �1O�0��<si,Nk�߃3�ܼ
�5G=B���]�j���(i�T$\��L��z�#P	�r�BG��C��[��V���<I���r��A�����\m1���0O|���_�|�M�k�� ?S/f��*]��#�aW!�۴)�ߡ������$6��d���J�{�]y	�-]㴔7�Z�'��H���rǡ�MŬ[���h������]`R�$һ�.b��8X;fwꀯ�j���߅�7p`~����K��=����0X�z����E� tN�rM���F"��e�y�EҶt����4���C3�	��i�a�zs�:�)��3�;#�m�������K#)�)���BR���D�R%�iP���O�p:na1��Zl�C�Mǫ߀�z��9R#�_;�i�����?h������r,[�ȳiJ~f�V��Wh8�5Ӗ|�Xq���>̥���E�1�����x5Rd�}u�x���L5?0m�L	�e�I�ԇ�5�x��9 �Q]dM��'��n��3��<
��D��q�"n�\��f����~[o����	�R f�KD���J���!���CɎ:wDs�(K��� Zu����3z�Q}��e�8�l.@� ���^3��֞@����9/^��<=��|K0.��\P����6��֖Q?3��W$
��S������'��ɝ�6[`n?%Y4W���I������~pCWN�~JU�&��X�IY��9�f|e�͜]�7m�߲zP�
�����+P��AXߘD�04���z������ࡰ��^�#X�b��5]Cת��w\�,���P�(g��օiϙP�i��u+�B�&����!�E_L��9�GʆғQߩ'�VXw�/� ����峩���Rq��njs��� IU���a�.h|�LB�܂������С�y%�I��z+�C���T�A͇�ћ�+&-d��@.$Y��ؠ'!�����n��-�`�Q �S*f��׆�q
��g_��v`�m+l��܊�G��0���V	�A����牼"�2NW�\lfä�=�?��v9��:+���p�e��d����sT��=L�u��
�y��2��~;�s^:h��I��,�La^�N��ђ�o�
W�fs�D�#�T�N��|M�D�(+n��ᥡp�8�}�sv��J\0A�> d�*+��^>qBND47Aߘ��蛑����h��"LLb���ſ$������!ى�J9����	�7ט[vO�:��ft�㵧ף�����0�[ӆZ�gZ�����n���ps�K_g�pP�#��G��.9,0AS���/S�s��,��/֥��r7�?��
8�U?�@h�`��rAΰ������NЄF�J�9����B{��nO���槠�Y
��B!���p&�(�uf>�n�)��	�%u#%��0�o,�&�����x�������+����zg��;u/4�x��$�/l���HY��"z5��jO�-�@����`�a�[g���U��F�9f���'�n��#���G�Gx��d^�_KH�ܲ
��x�t�OSjI�j�{�}�~��d���ȫ�4���gHl�!��Xg�����Hi7Q$�M��K��/��Q�6�5z��a���GyQ:&�>>he�u��L�Z� ��7@�	P�vI�VGﶄ��tt�e�a�Ӝ��6����X��6�|���ه���ޒg��ge��H��&+Q��@���D֋�(ҽ�F+x��7�c�Qzӄ��\ge/�@��P������z���Q$j�>x(U��P���lAK��`C�}/����~9?�P�Q��H_b��&�����=�)s�Š�A%2	�ƈ���z3ugz��I���j��7�J���Z�̩z�Wd�Z(�b,���Z�g�u���r~�at����c��!�h��.��/�k�����
��f�x*��i0�"+�YiJ�v<u�DQ�їx�.n[�������.	�RN�|���`?kru��s��ϔ̩z~R�=Ьt�̖qq�j��u��꓄���#7�f%��������}r��pk��v�Hm9�_��Ѥ�z��������G��:�~�!�<E<h�Dol[���uqUk��[1���������[���o�Ңcj�P9�[ɝ"�D�\1qAP�ȫ��e�kL��d�����[�a[����US%�����t������c�k�桻��]!��4dxS�
�d����q�&0�FRUٍ����i'm}���"_�鏊`V��q�a�r��^g5'f}|�/`[��?�l=����$bA8�j�WR��П#�(��!":o�緃�,Y���`@�8�(�4��luM�HqZV�r�
����B����a�;R��~�Zd�.i���=�����v�NP#��sz���J�O�J������lሏf`q�'�2�)��6�d�hpҞJ��m�EBL��y`he���χ��J���dR�m����hɖ��+0�Tz��[Z#B�&[��:eQ��|B��DA	Bұ�]'Wk� U �����u����X�튙���Ao�D�� #bI���|Uz��p���}yR���MҀ�@�%�[����%n~�bB�y��[�l���Fi����Qڑ����&[BQ��B���_�Ҽ��C'�ޘ.�aB�ZZQ_ZC4��^�7�4+�r0F9�p�K*�)&Z>���
>t�}�����񢥊«�/��鱗۱��T�117R�1�@v,tUu���%qZ�r8��[�*��_������o�q�^Z}��R.�n����T7GQ�U�m".*rv��m���C"��c��*L�>Z����4x�)a�ޖ����r����,
z��-:_J�����e~5��D�Չ�_����J�x$Æ�ʘ�;�j�ˈ]�����8�8l{��=���@�l�(&`B��m���v��Y<<�!f���)�Kew^�7����V��q�$ٞ^��C�GtsZ/6�Z��C�&`�?�ur�v���>F��%��v*�يu�[H���Ґ�^2�/ƅ�4w�d��>T)��b�e Z�"��	&t��,�1�HL�ȃ���A!�B� �y(�R4v)j�0�В�L5Ħ��P���d���q;�͕�2����eud'W�5^TP�^dxfϵr��|����d*;a�:,�IMM�f�q��Ѹ�u���Pn/z�"0�f�*�������|���-v�=q�D:"c���3me��v�F ~�Ԯ[T>����|q��t�sQ�#�jE�����$x����vϵ_[�,l��:���t��Q�K��-
J���7�^��� ]�S�� ��:��"�t�^�<�%����e���V�:l�δGm ����,��G׷LJy�rH�,5~���b@v��Q#�I�	D��7�>�h1�#�eMe�����TY��=U��I��I�.��>����0�N�@e8;k���R�� ?�����k�dfr؜ڌ�����Q�j5;�>�eg��us\�Mt-\.�;8T�ԃ��N瑝BᰰC�ٓ�����}ɷK��^y�����p�tQ�L���w-����Y�;������zou5C�Io�}����+�s���0�(���t��:����Fk/o0���&�EbnoQ�¢32��T���������x����Q����l�,����R7nt|n���L�@�P��o@�G����BfK�x&$*�*=�Ʈ���=p=��󒥄���;���aT`r�UǤ�2�ѽ0U<��]����h���7�o݀���kK� /����EŴUW��X� ��[,Q�V�1y:z��WJ�Wl�_��������T_�]�Nn����[^B3fR�lup�3,�$��&v�����oN� �G�eߢ�FS�~;��2I�+�A�/J#xg���(s�<�G��(8�Z��\1��Rԩ�S��qi���u��x�$�.a���[>����P���̓�!����f�ܶ��)�(�����o�D"˳p����S;���y,���4�W}�4v4�H�.I��k ���@7�$�"��u�k��.V�> 4_��\t�:^)��)�~��b�P$F��u�
eͱci2{[���6a}��5�(?uLN%Tr�Qb��O��2-I]��.8�2.|�t�aa�E�/��K�P8�h�7�nq�8��AA���XlxVHYEB    fa00    1e20�|s�2�[y��\h���$� 5HUWW��n�' ;�@�Ԇy�V9�\��ȸ	}��#�x�Nô"�y�1/� �~l���$rҢ���ύ�R����k�� D�n�����x�U��0�Z��M:̈��O��}�*X����xkx7�o��m��@f��*���|G\ے.>`Ś������4I�,mY�c��&-~C� �՜�D���f7�e�r��d�q�GQ�8��J��)�+�Wg�]�����c���؃�%h:.��"�X׹0����d���"6o��2� ����WY��=�B�x����P�>��䇫�)��û�%��Κ�YE!@:#�K��3���k4#�K��~�4e�zݟ�Q,�� *|C~7UzmK���w�1AI*�ʫ��(�bcI��mQ޶��������IQ�'��[Z�sIJ�|p;���k��9M����Od$n!��ř�x/br�JE�Q�Ԩ�W�׊���>L�z��S6V���m6�v��ό�˨��{Ap{��	�n�p����"&vg3_2y����gq�5��n�H��(�ˀ~�����^V2p��q�j4Y������(���	�����;[Bz�G��F�gHOpްb�<w���_�z���
���>���rX,�QP�k0{��Ȭ�Z�O.u#�bwU�X�6�C͐���߮�� \�����R�����/��&�_��?��|�K����ʨJ��\�!��Z��C\E��|>����zC~����GO"��pP��qϗ}O5\��d�"g-��^���:;J��� �����0����,a�#t�eis�z?;����k��Y]�[������?$�|��b�R^2�W�b��|�ķ�ˉ��t@2��F��q&��*t8)p'�m�/He^� 7|vn�%{+�i`�A�ơ]Z�e`|l'�-���w{
c�\�� ,-���	6s���et���b�G ��eLq�K����7op��P�W1��%,tl6�\��)���7�n�;E����Y�p1X�	ߥc6�ѿ���z�i��i�R�9�	�z]࡜nQ-����R�YG�����tN����F�2��.&��yU����`l6�Pv�=׃����4�����/���qm�i�i.f�mb����`���D�������}I��"o@�$��B�ֽ�V�Ո͝�c��
��ՠ��&0h�4%`n2��GfL�rڃ*��c��!����,R��_�ܴ�(�vCCB'�]y�d�'�_�_�D�G��g;F)Ql�j�a��D��+��zQ]�;�o����y�`�9�}����D:
��e�7.f6�Ny㿉�{��U(B���`����ge���ث~��X*�j 2��MRW� �оt�Ui8F	1 4���z����������H�?�O��/{�E����	�6�Y,3�DeZ��3.C�{	����iST���h1�'CQd`pI2�uސ��5�^��&H�[��6���}`���ĒZ��;U��Qq�"H
ā�hB��L�W���J�@��+�������"*aR/�ް�9����<��8T|�o�"�6�_i��a/�T�5]?���C�>i��^L)�Z�Zvi�:�61��iCH?������5#�7"w�(����O���QVy��2���<�?�{�������8[���Li1�slp�z\!�}��o
��*A�\�^��]_�r������6��c,��N��c��~��`�����r#�E͸.D
�\�������g�̑ny�	�P#�ޅZp��)���Pb�;yv�z*�m��L<�8/3@:��ȟ�w�K]�G��ZOsl2݄�^��P�a�pm���!���(8�%��Y�"�f���[(���B�E��u5^����%�V�-��;���'m��X��Pʆ�9�^���^L��5O4.H�;O*=�.4s���'#ԥ�U0��r0:��L6�?;� 	��&���=u�_s�|�D�|+;aS��6Ϻ���y0��x�3����{_�8iɧd�zT׍9Z���U����g&ն�W(W�9���LSL��	���q��Ι�Yt��C~�C��DF��[�ęGAvϬ���[���u��ln���i���^&��|`Ay0l�XN8���I,�#	��S�6(���&�,�r��o�N I��[�����uck+i����P�� 6�8)2� ���*�MAVDn"�T�i#Y�V[k��CKs��99��f�:;k�A2��]�lA\h!Ia�@��ٴ�
T'��N��D�
|\�(!�-�Y�SɊLeՓ�/��j��#�8,���&�2�x�§kWC�'Vt[�>m
�8Q��� |Vk�M���ؕ�RH�8��]��vT���Rmg6{����4����������D/a��|�}`|\~��8�H�ou���^��o���Y��״]:2��!t,�/^U�%�B����u�y��פ�6��}��خ�����-�g���x�V�(����p�������[�>#&Fp!5�NE��Gt����+��aZ-��|!II�=��ǔTHk�3���& ���������n�������	ܒР�k�O�?��B8��?3�� ��+���P�0R"0`�@�������U��{����_:�C���0�1R�+'��D� *D�!mu�Sv�3쾩��{�l
Th�pcfq:C���/`j|��W]��
V��YZ�a��SC��ft�F�����T��{T�;'���dRq,������g�|o���Ό������o����	}�ޝC!�JOwk\���΢Y�]�#�������K�F��x�9C��S�	�����Xԣ��dԓ���ߝLu�
��d/���'�%�L�g�%�Zk/�B����j|����f�!6ΰ�(�� sHc���Ģ����?�֙{��gG�I�q�G���SA���~V �`�,^=`�=���	�M !Hfn���[����P4/�&썘O(&�+k�����6.�-w��,�Io㪫�e}_��L�������[/#���jJ�F$��:�S����If���wO����h�>ߧ� ��HR��F�Њ8X8h-�e87_j"���@���!yh��W�]�?�\�uj/�ߧ�8P���G;�" aGb!��KL���KP�(��|6��R�ddx���>�����=��P`�p�n"�EOxS�[m9�&[���x�e��־�
2H$q��"����&��j��J����l(�\�Y�3	��b��f�~3G���_�^�e�y7��3;���M�wx,�ܷ9Q���#��i�/uB'��L�X�9�,�ǂC�bHň�C�C����"ʟ�<��w�~8Z�3:x�IkG���$��f�4�wZ�٦�Ɛ���4М�d5����d��1B��p�cY�	˸G�I"�v�3��|;19��%�2���0�����)s��0oﭜ�=!v�!��W�Js�В$�On��H���(�V�VC��*;ޔ
q�	m	�,m�Ej`�F$G�e�k�4�����J/��
�dM�k����7��ޞA�C���=�R]Ab��ˏ@�w�&����8�n0�lK�Hn���t� _��[�\,��5��+����Ǩ��ں���Z����5�/+Uu�Fk���^���t����pM��P�+��@ǖ�^�P���SO����~��ː�[+��٬�Wtg�������e���E�$���xs��]�AcB�~��^rKУL�O�8B~�u��?��&.BK�Ə�t�p$N
��tR���x�6���R?T6�cf����鐋 �E��P(�Y��J����0���6~���N*��XE?�e�!�����r�x!#μ��A����w?�v�O��b��E�ej�m�X&x$li���%�{Ϭ
��ם�ܥb�n�HhlE�!�f]W�Az�NC�rQ�iQ�\�K̸'d�XIE��e��G�;��o��!�9�MW�_�A�a��U�`=����_˔�	?]��s����z��ap~��l�6����������$_�l8c��Z:��:��t��+S�.V�i��*���|�vp=��(F�&�E�U���}\6�_FS���'�W��x�0�h����f�Rm'�,M��'M����<�b��}���Jfj;h�Pv���)>������!8���k�b�'��b)�&�S�7`�pozR4�se��|�(�l�
Q�Ojb�� rB��Z�`O���!��p-U����M�-��_�B4��W�l�x���Za�O��5N�f�Û�Zz����5M9�l�3�=VNHU8�P�#��itD6��.(A�J:���s(�ͽR�!j ��լ+�gLr�Ʌ�[�:�4�B�&&���V��x
�p�(��Fm��pp�E�'�f~Ï��K(P1��z�~���Q��Lo��QG~ՈR�#���N�bQ�N�挮�M<�|��Vj��p�A:j'��%�o�������e6� �6P{LvA��5�0vË��>w��q�(˻��!�H��"e�7<�l��)���e����pp㻏��Z/�1�d��kn�u���j�2Ό4��`5��t{6bs4�gJ���C#�:*dat9.Rs�Bj#����
RyL�?��/��Ў���ʡ &Pl���H�E�j �|X�kW!�j�1Ut�aZ�q�@�/��\���Tёr�C��8J�L>�͞�|QMT>��5��<Hf��k�|;���|�ɋ�dc�h5@�p"����_��q��h`ad�w��a�1���J���ʂH[�ƳP������ S��l��Y(C��A2\˱m��nbQ�4�=Wr��S��+#��n�?��6�[æm͐�C�+0Ƿ�3���?�q �@�'Z�o��-WR�~�[�Dv�H�FԂ�T�x��wE���U��(L��B�5$��|[�V*��_�9<%� BIL��'X���W�?���\��=�A�Z�v`V��+o9�E~��[�� ֌�fDL�#b)>S�6;�]�"s~�~�'bp�����%������*�#�X��o�8	!)�<�h�Ě#��H���1��&IL�e���
��n���h�t��(�<�����)S��|p��=���`l�E��/��Ŕ�;k���%���%jU_�������oƊj%�����q6ek�F0�M��X:m+��c`y�<�bWR��>��`�~C{����{���VUM����Sp�j6rE���W�
� ���-"dl	�z�o�4���h�=�ڲX�3�]�FgAC;����rR35aj���=�?O���X�h�_l�0�m���b�|���R`~��~6��)���M�޼܇�V ��Fk.��w��\L��-���n��K��ժc$fa�i\��G4��91:���n��.F/2�����N�
�P6�	RjW�. xs������b�8��&�����u�S��b���i�*�?C)���QѲ�N�_��w�+�J�s�\��F�Q�U{ ���j�� �QX�㧨���<Y��W<�aU�#��Hi������ÅLb͔�o�,�=��ph��뚊���*��)!�~�&5�e�"�����#�3��f|nlj��IY)#x�>�h� f~�C�-�� ��pt0��Rq����L���⣒t,�kI5�̧`3�q��?�q�o�����0^8�
���P�fj|��yV����v�/C>��`�]A:����4�ֆ�2U�t=߄� o�nE{����G;&YL�j~P1'�^{���1N�c��(@E�AxUog������n�z�����~_���òu�A��`��b�35QdasN���[��YU���3��n��d�Bu1���q\:ך��ݴ�^��>�$�S!V\G(S��U:��6Uvuy8/R(�C�-b��s�Ӯ�v{����vW����r��������b-q��&ֵ���m����V3z4��]�ԝ\��:b�뾌%�A�d��C� Q�8��@�s�PV+��;����C�en�ҍ� �T�!��F���e�a��9f
��t������-�-�y��I�3^��4��3�D6�[�{e�'�D�=H=9���8��V� �P���v��T� ��N?^������+F��9�"���?��j�/�����{���,m!��ۊ�١.����,��P�i���=x˚�[ZAmcr����3����ś�Q�-2&~s���g�'�Y�����+��=�������c����U��?���5��:Yc?y@� r���2:4���B�A����spmk!/G�J�`⌄&r"i7� c��_Nv�
}4�CZ/���@�џ.�`B������w\f�NTϓ_)(����.>@<e��Q����!X4���X�-�;���E0RW{�3�s
�~C����r�Ϭ�2B�u��"j*Pw;1�1�j�ep���{Ҁ��K������X�ջ3�|0�ݦ���|�o]�g��Y-<u;p'������mk�U&)���)!77���g�2^�֞��D��9�0L�?����\0RR �'�,�G7u����k���4(jP����I���n0 *���Dr������HI���b���⌌��� � �2K&�y<�w$�i�k��kݤ�m���*�MmX�z�������fq�#�sMl6���K7nW����L{L��c�:�������`��pr�<�o���(�$	+Gb�rʍ��B!`��3��T�v	�Iݝ�̋��� (f��7�FU{��Sql�,�Qu�Fàp}�ݎw��[^��א{e��s�:G�>~��.'Ԁq�-mI��w*�����V{�g�	y&i1�����>%����'+�ni�RG0{d-��5��\�*���ȸc���)_�$���0p^�T���w�<��}�h�t�g��K帛��ӓn^+�>o�TD,�bȥ�J��������z.�U��v0Q�P���)87���W���f`B���n�#SB_�wsH��b�ś�w&��Si$���F�.��9�@2��!ıh,�䋩(�v9�"��-*�\j^��к-��|H�]7��4~�w��-I�ǀk0���I}&���1�f'D<��D��_O���&���?jW<�)��	�����eO�I�_Zނ�(��:y���rE�&N8�����Xg��^q�8���f{�;�7[���xv��"�Ԭ��^"�"�#�%�\�d��9�0�fOs�Oj������d{�������ef�����f�L]�� :nRAiW��f�7��ǻ�����?���`�7�'��m��J�L��{b_n>�5ޕ�q�:���Le��,Ǹ��!���4��;��J��)[�������%d�bBʇ��ցg�QҼ�ok��~|9����t��x:�f`�a�����`�C��Lەѡ���ɲ(�M#�"+�v؇��df���Js��ů�	�WW��9Y��ا�8nʁ���%~�&�v�K�0K�g ^�����XlxVHYEB    fa00    1e50��햿�&�s�iB[�����T�<���)\��)q���7+
V��sԂ��"v{�7�s�����C����$�\RϮ9�%�A>��׸⼶v
W���!xr;b�d��ܬ�gt�~�t_}s�1���L]�Z�`�̒� ��Z9Z@2�/���}��vH�8�(,�]�q��=�7 ZV� �X[ħZ�%�yƕ��OP�;`!�.Ɛd����
���_��k����$���Vq�Ir�Ԇ�B�Cx�yqN��0����+�})p>G���9���X�̽�ڭWep�s��%�p5�S�?��<=d�)2AUiZcW�������g���]p��(t����M���]�~���zh����u�V�}&u�p�Y�@\`�l����ڞЎ1���Fnks* dca��+)�cE�ď�+
a�h��kY3@om���ܫ�/��e2�-�5g����0�"�	�Z}�ž_��+�L�������Vn,��|Ҷ��>?�{�mL���F��@��������I�����KA⽙`6�6��-�Xc��� ���C�C�m��hL]v�؏�@�Z�4K�VX�f6��o���'����K�D���B<]��H��I�A�d� 爺��=ʤ����HV�S0������4�|���������L��:h�t��f�1~V�g�bdA��Y%u��8�ii�����@.�Z�TػO#�.S��C��;���w�1zz�����
�h?o��]]5��-�$���~���騼ɶF���
;���čW��PPoI+a	��XCޤr�O����,�i5A��fZ�
Wƪ���2G~3ϧO��ֈ�^@�d��
ˑ�S�
Uc |VS�W~���)t�E�ή'*�N��xb&VM�lb�*x���#�v�'	;�7vMWFa��Ō�#F��`x�9���\���p+���!� ������V�9i"?���&��Ĩ ���/�m@�)P�,�r���V�%��`-�W�`�(�h�;����J�f�T��)�ZH]S=�r�(���!�����K��'�0mЩ�����e�9��cL�s�@p9�W�#��f��}U��{ ��א��D�����;h�:slE˫�i|�Q�d���`��F.�sΞA$jE�ն�����κrfnh�=�[����i�)���"oߍִ_��q�����qe�����2�[�h��Hq��DXc�0��O�EBd�h�?V�����]����sl1ň�P��\��Ԉ�N�?�6ęv� ����@��O��X���J\u��Qs�~a]y������/ȷ~�Y�"�E'�[?-�}�:8/��7��ߦ"�q&?9W�r��	z�AҐ��U�[�.;Qk�y�B�+hܷlvEu������`.j���,�����7шba��M�A.��
o# ����E��^�m�5\-::������{>'�gS������e��[41H�!?�@x�;	���2|$���Ml��<	Zm����X����|��H�6 �$�}�_��(*��E��s�����������a��2|�O�f2\J����B��b�w��oO���=l�b=4Lہ��6H���k�-6v����O�z���藸��J��(#������-=�Q1�LZf[��j���L�XQD<n���JE���a�*��s�@ .3�'��ƝL	��v���(�i�O�oHŢ�����p�O�W���J��%�����)�B5���Uk�Y8y���I?���}��Nm�����Qq3%l�O�F[G�Vn}�$h��I���_�&>:�����3���*��]t�sS�����4�Ͽ�G�0��o�W RϦ)|4�7�c�9k�>�D �G�#�͉��v�=X���<���;JKV��2���Ґ�x��=`ޅ�;=�A�b�Ri4���u�;O�"����Ug��`��0UO�̷^ ����Z|J��Ҍ� ���6Pew��Lu�h0wz9�\�Ϛ͕"���E$�K�^CQ���x�	� ��t�Ix�'��l�01�����1����âYZ"~eds�2�S(忶�`�t��r"0�{$��8�S�<K-_#p�����Lͧ�h���x�-Y�ܭHL�ޭ�>>�Es�8mE�t`'�<Ke�@ p
n�8<�->ek}�VP���O�<2��
Vr�����Ig JQ��K��`�^��\��zJ�?(y�+��b?*:�#���\*�!,N(#x��m,�ߝ����'�����dCuB�Y��\�NF�[�iX��Z��A�^@��I�.�H���[�T|V�9����$��*VΜ#9�}�����Μc�@J}�U���P�)�y z�i3�젘i�F�.�bÀ=�d5ȹ/�i����W�?��zk*��U��I�n�;��Y�.-�Z��>{É�E�`��-�y�^,�6ec�����t6_��4�d�C!�|���z�6��<=�m�w�.=�M>~̭a��J��_(>�ʷ�O�� {��fE�n�I�M3�>��R��*����RW�>_����*�R?���<&�_��mO��#��\�Oz㊽��#�Z�w�E�CXF�����ӪuV��?��o:d��B.ˉn���2���Y�b��ՙ��?�Aʳ(%.����ޟ�Q���z̮���>�i�ׄ�i_�Β@���΃�.K|d�q%��,RwK@���B�[1%?���FQT�w\���5Ú��>���%���G_$ڭL=�ir}Lj�耟'�G�	�1"��m^���o����;ǽm֪U��.�?��{�t��`G�~b�R���J��S�\�>�$�
Ã'&j�8�O|�v�O��5�Ýs���R����)Ӎ�)���1��s��:�G�"$��c��',;���9��az-L�Ρ������I�H�'�̃eͻ0u�ؙK�Y<�U�69Dq)i&� g�3�_��¿
� ���?<��Vvd�b�vEǓ�M�X�$�u������NSDc�?	�hGs\��TXo6b���0�{� ��?�6�[F�Y�u��069n��"���Q>��4ts�׿/�t~�����BD�ڛ��@��	�#[0����b6iA+�V.��c��v��6���U�G��h�أ��ټ� �/�g����scbL��-��e��@v��󐯒�zfz�5N��J�i׈��V&��y�5`��$�g�,J�+8"c�7��k�)g��d�ɶ҃\��R�D^/$A��NPg�����{�`�Iw��A�gs꙲+�sR���3;2�V��5�#�7�Z4ձ������?+��d��}J��n?"P-�sO�ف:uvCba��{�@)��TC�^	l�r7�мL�햬,�N���5�{���\D�4���0\+Lis����Eh��-L�5Կ���6F"g%dN���o��KI������F��u^����%�	��ҘX�L�35�{�-0>�)���A��\nĿ<��]�AUbK#�Z��)�p���&�j���do����!��~�[���hv$t��y�zA،���ɍ�C�;��/yb�_Y��`#�m��z�dON��uŧ�Dc�K�B�K�H�Fcu��qS0*���z�#٣�ە�
��ߟ�>jQE�B(�����
�}�y�z�槜b�N�4I�2ఞ
�V(7`�����s=ڳ@����/��U�b^�ޯ,��vDA9�uaqa^���1�N��(�?%p�� @��y�ۓkH�������ö�}���A�CM��2�ն����	�:Ԭ<J)���Ab�-'�,Z�cᦳ����7�k>B�E�kԭoX:::n^�ĸ����7XS�ؒ��ɜ���)��/����E�s~)�~{	�R=߃ր�6BB��7hOc�Ve�Y\ԓ�m�,���
�JW%Ra��|��ӝ�=��_��1[��듣�g���<U�lp�������fUOX��5.���~?l]���l]��{K�?���@���$z��~�Y�?�!K���3��!P�����#V�(G�g+)��G:���$@݊���P�8�tp=���̆'���o��vE3���W]n�Qwe��T����.���l�[ ��x�Mh�}�u�#���W�s=��T�*��$斣E��z��~m$t�'��|��x]�М��OS�ݴL1�YcS���G#�5-&��R"�|�CX���pe��(�Ur����:���2�~:D�	��*���W�\��L��=ᑄ���j`,��, 5�oduE���@��3�fu40���^\v��)��l]������h7�!��+{��3�`�J^�'���#ϐ��1�}�:Tz ҭ˽�3�  o,�@�`yx{L|C�f7,x��ď�z��? �bu�5H����:HE�w&�1$D����
5�L�R�,N�e�}�����#�?�/$�a0y9k��3�
hu��,˙mK��f��;�~q�ːFfF`�ÈE{(�w��
�M'OR���:|ٵ)�U�Zx������c��a�?���yk��0�1����,n��������
2o�SVD #l��B5kY�a,�{w��BH�y$�w��2�L���R���HJe�j�(/?�*��*%�r9N�_	��!��.�%?�o�m̧%=���H������N�}���z���1�A��6/��N��"
��Db�����<I� �29����*8Y�̋���huQ)M96����!6|���CA�o��`h���-T���Q��c)7#��SSP��N`���_�0=@(�屢� ��;��|r��O�M#��--]C]�o��Q�Ε��
3�*ɻ*s�ܩ���F�azV�
��[*+xQ�z�Z��V�
b���3 &w��N���a��'��G��U��/M+�9N�����^��hާR1y�j.������k/r���/�u p�r�Ɣ��*�R���L m����Z]�{��������^#`��.$K<<!hvU;���r����u����^�|���/}��G����g2Eq� Q2��R[���[��F�����	�����Q��]L�o���v0��*��p�Y�u��q���>��ҶToS�2)4âY/�yg�p�Wm�o�7��#����d|b6�d�{~�"]Xulj?T;5�m! ���,,�ll㑥��~��Mײ����v���ۺ�O��}5{�.%�4a�:�Y ��n�����IQM���p)�êL�4�RD��fE�S~�':�>I���.z ��X�8����u&,������ѝ:B���m˛z����&DrӼ7ok���̱���7F��z�@5K����=p��o�$ع�u����0�uD̼��,�wݖ�^�{�&U��o��$<������k��B�MW���3U����wM7�H(IyM�㎹�拰ݲZ���דg��]�T�u-"  ��P�KچY����{Yp.D};���v3�l�:J��>����ڣ�%B�7�z��kk3x���[c��,��}�M�@�Fm�ig�Đ�����Bp��Tܾ��&�V�ﾒ\���&L��p�
�/U�Mv�SE��!r*�	�C��N��&���'�(���}���q4I����\���	�6$�(���-����dor�.	��M`�\YT��l��p��Z9>=�v��щ�C��Kh���-.��n�Go�kd�p;�"v���_��օ;B#*�V	X8c���ˮd�O:�m ?��}L���*����g����wل�몌��C�C�Ra�-��q��?�fݧg4��O�Tq�1�n�(�)�2- �l.�u[��m���.Tyۍ��z�@�oOa{����������n0����Թ���� Uٵm��Mh�!�w^��n�I#*ij��p�%�	�0�a�O6L�*<8�^N0�C���c%��mv�+�US��_$@,V~��(ց��_f �
[娺�ə�
i0�<�������aM%�[Ou!b����JH�̙�V �@Bs���k�P��$0�'~�u�6�.s>���N��>p������0���Njڰ��G{�Ia��V:�r峅|�b��1��s�q�[2՛��6�?�K�� T� ��'�}`��pw�	y��>�Z�Cd�`u�1�8.|oP\�L�[F����5W�mo}�33�;�%���p��'Ju��t��Y��� `d�C*�ݥK�41��NFP����]�hqǕ�[��1�}j�jnƁ�L���Z[�/��߬����֡̕S�J�&צ��QZ�*),O� �ܬ��$Za%�}S��h��>�(5��T�aM�W���H���l�n}N(B�mt�"��ᨠ����ӌ`0��1gZ��qA�b��
ݰ% ��Nh�8t�O�+�2�oV+��G�:��C5i�@��`��e	���Ӡހ����n�11���x������If��t_�	2�a�=ńPxYi�}.��D�!~��a���˳Зv;��ﰿ�;,��x'g����r¶M8-�'���!��bN
��o�>1�L�h���y�Grd_����i��&��������FB���2��O4q���ؗ�W��K�JA�o#�#�T�z�O�j:�<cќǄ�Iq�a��J1[7�i�ZXs�3FB�|����6a�{\|U��L�XR�L���D�b���.�A,�޼�A�?BR]�U\0>���c�a��Bw!3G �L/�O��
��)n��5�ۤc�^}��Ti�=.���ޤd�a�{��h����W�wX�SS����>�4�\-���}֤�Ȼ;��[�*�o��Kz�ނ�<v�b�_m��Q�y���pq�7�F�b\<�ILH2�:��0o���2��]3_�u��8]9-rd]iY��|�m��
Գj�AW��HD�v<QI�c<ɝo�-�\1X����U����s~v���gmP7/f�ڠ�C��H�ORY�."�;���`�~hA=�0��c$�(������S.��gz�']R6p�M��������:�B�y��d�Tˢ?�!>#�C�*���
uH���n �܀W3@�_~+�d���H����.�(b�~��	0}��&sJ��y��zW����M����Siq>��U�Q���"4}5[�S�� +�]<Ա��ɟ��;1�����O��{�z8׵����p�yJ��_'��"�G��	q¹S��%���ݘ��J�-�ǋFW�����������/NE�
%q�
jF���Zy9t�����
�p�vc�Ņ�wr.�� T�=4Gޚ�0���y�K^�ӿ�Z���c��N�g�ݢ8�C�%�P�2�V��0Wгn&䑿���_�8�e�[D� ��]y���&̄�Y�H�)�J�ߩ��4E�-ɉ5���?���E%�88>[#~a'�^a�7BEV?85���2���w�4�R�uy*�=B_{�/r8���K�yp�sV����Ѹ�M���!+�=`:�i ܲ�������`w]��x���kk�s�D���G��Qt���)l$���Z�����2������|(�8�a����"��J��&��4ԸL��.��;��,3Q��$<����cӔ��-D)3�x�U��L&��].��`JY�{���B�!˝��>���BP���%RM�6iS����1e��V��(51��I�XlxVHYEB    fa00    1da0�7��ذd���U�����'��"����f���N�2Q1a�Z�dZ�qw��Lv�c��l���h��o�,��,�\�=H�3I�q�E������%6V�kD�"�@nŴ��oc��C��CތB	nA(�un8�����Ԏg�1R#kb4��I�	��P5�$}� /�1��Uj�{+���eCsf�X�<_�H��XEl!P����3^�{��re�����]Kܧ�Z���pﴹ�:��	C�CUț��L��Ҡ�������	S�u�d�3�HZ���� :g�j1��s^����_�dt,OI3ڈۑA�
�����32�O$��%�;���֎���+������}���#F��x�R��+i{�*�|�p����&}id�j?�W��Ud�PA���a��xVo�qp����v�����#�i��MNu���@��!��9j�ȧ�u��C�s΂���B���R�������|�/W"��� IZ��XG�Ѫ^�z�x"�:E⡢ZBW)�(���C+6U�EƗ��:ҺmZ�Y=��%"����MZ�)ǭ�l�Ö�RѢ~/e�I�OPn��z�Q��d��hu�ߜo��i�cs����W0N�;a|�����4Ns���JB���*+�! i���VO��1�h!p���C f]��bH����A�GZvb<����ŕ�9\��s.��	 Ny��x�3���_�:����cc�$�����a���B�Btל3v�.���HT،I�s�:�R�� n�UṴ�>��Z���w)��d}T��鬀4'�H���1��� Md�[����Q,Z��'~؅�;�$%�v�6��Gf�ğ�r[K�T���AlP!�lKl�5�!�V��?Uݮ��
P����u�GZ���(�N�Ő�|0�lQ��
UQ7E8����$�m��n����gY��/����
dc���&�@�:�\�ڇ�1�=�T���`~�g ���bǐ�_�����{�8oNH����-'ʈ}&�����%%��"�:��5��������y��l2�ް{EBE��h��ũQ]L���A�X�u�{�����Ta�$��Ov��,�<y��ۯ���v��	���㽔ԋyg���hF�5�.r���,M����Fj3�<t��G@�8�sv�
Q��R��C��*��,b���Dc�?�N������]�����*v�켴������ט���D�ڣ3{!��un��tR��;�+H���֭D<��	w�'iKbz�fZ�9{�����:�+C������2(}N�Շ�V�U8�>�5�*���m�P1��4��L��(�-�S��R�VL�����2ɐO��Z.+fYD��9��5^��6�B�]��ŷ�j�`W�
[�L2Vҿ��钾�{�ⱜ��ik�ZƆ� ғo�f�v,��]�/T�fOs�?�����1�L�9	4�''��ie�οɘ�u�8��5b?2�"J;C$��<|�<�����(����sp��n߽-�dB�`.N�*Az�t��ǃ��ypx���9{��M���<�bZ�Sp���1�}aM�g,���P��̻�/�^� ߤ�?��J�^"��l���_D���`�l+�������0��ɀ�1@K�{�.�?��j6���i(�F���8��\\���1d�[[R��
�_�"����xTe~ ��	<;Q@��4X��e!q��C�*R���?`���F�`�!��e����p�h�P�u���U�!�v�c)��a�M*�8y� A��UKsi(T��?����D�k��4�)���$>w����!zU:�2������!������v̸^G`���z��NY�8An�8���y%�����؜R��m������F����%TQ���5�@��j���F�5
�&�)�ۆ��<�����@.>%X�V�
8</�B)q2��K��6 6���]���S�oJ��f�aqx�VK��YP�1�Q,7�J��$�[D���d7��i��� �1�`V����}
�� A�XA��&���lF\��+V��]�Q.aJ�f�C�2�������6�_l�,L��a���a�
J� �lB��eP~W�޳E�?�+s���.3q/MuZϔS���u�*m�D
����2ѼD��+W,��F
���k+�)P�;����9�-)��^��!����/L�.�Ow,3�-�&+m�C����b���#��o]@�O��$�m	ʽ1�X�����<F��ǅJy��4;Fx�r�^��S-گ�����Αن<�iO�k&�(u��Gİ�{������4<�\M;)�����:���}�_:7BS�aO�9�^h��nr���ˤGH�ĒTh�AhR����f���FU0D\d2w(Zl�E�(q�����k"�*`M?�9��wx_�fQ�I\J�Ȗ	�臣������iZ� ƯP*H\�;�ϞU��%a�^�q�*)�)���E�b�0�?�]9�(Q�E��<��dɼ��s���)R�K#P�#V�H�g�g��]فC���N5K4Я�l3*�y�W��Lᙆ=����oPy��W>�<��+ɛ����W��Ӹ^���ج���)�!��9��\�N��~k�S�'�Ā�Ã���m��㔲���kŐE�u@ƻ�R� ���O�;^; ro������G�߲^O��3�G�RR��1�м���1(T��e�{ߕ����t_�U?��h���ݮx	NJ�����t�hZUY������D���w��`�vV�]��]�ˬ/��֤���wwX�9��|�6���2Xgi:��B|�$Eb�xJ���;{G��*��.Ք��Ye�ȳ+8zċ|Z%������h���p�k�hPi�&x���]�е?
�ڥ�vs������uQ�k�I����bB�!5)5ո�CK&�,kI�o�;�Q-��)�Mh�*2���QF�ɸI�`� L"�?��_�0��k>�˨����s�J��ƍ+��Y���ח�30�1�[�^ }�� �����CX��2��+R�g	�>@����٬)�a��~���Z{����"~��W���G�]1�D�e�,Z�z6��� ��ʢ��waG7e�yh>y2},��6��@��N3���|5ؑ���'$O��Q�.9:��o�yr�����y�S�J���CS�)$��+�qj��m�nqw�ma���wĊ[I����rU?OE}������}��)"���U
��EF�r���B�����#��T{҈�Ӡ&�t;š���[�|y�tY�0�pç�.����B�O��U3��ΉQy9���%��^�8��Fs+��|$dװ	����s�"�?P�.f��q
|Uq��q���~[����s�x�k�b:d;���"%+.���t>�� �$����!O���Ȋ���{-8�G�"@�S�!�n`xV�o�&`�}i#&��#۶Ra(?l2��-/�:�Wv�$R�ak0�q�p��a���$��vL���?����c8�����F���]}���,!�cp�5���$�ߠ��l��447�a[����_,���{ߖTP!h"�aj3iύ,-�ʴ��(�tT�̜�B%�M|��t�Ɩ(��t�wZ�#�z{*��L������+���B�^�̏�Z�/'F�����]������`�P�@�5|!���y�K�6����9In�n��2�� -?,yPo�^����mR��s%�v5Jh��d�/O]|���������C���W��b�	W)2��3�$����K1��AE�F8�9�������o�5��ř��t<�DE���P�ПHɊs�v�H�e8lڽ�Cj4�yE{�v�1��w�2����67n��~W/A�M�2��X^B�<G<^JB�d���&Y樂z̲�N�\e��{;��y+ZO��N+�j��������:���1��� �7�����&�?���l��	�q[�z�J"rn���:�r$��?=f?����'��=�=�d'.�m\5��$�^�hȟ�O��Ž����Ӵ���QxfhTb�n��][��xp������Wy�\o�AMl�6r♎���P7���e|rUW�2<0���󑪼��:
KƎ�p�4��� Lp����������l��� >�����@6�ۤ���y�����J}�P��pWt���b�{�K�ie����Hn� ���k���?3��
����8�<���SSl��~�!��|����j�X��)�T�4MN���d�w_��[EÓ��P���euh��F�Y݂;
�O������M� �:X(!o�5�O��]'���!�h�7.S�� �	�M7�r�yoW�)mv�u��&�YQ�d&���Ύ�I8D;ra�t���!�C�i_��������^�ˤ@jid�<9"ᝐ�t6(��F����.���k ��UL�%4龤Rn����J6^7Š*i�|Q�"�,�_�N�O�}��_S��¦g1�o�(�{����t�N�?%ȭ2Հ����N������K�6�w��-�&��M3�q���	o�CȲe�X�K=L�`�>�ex/��=���edZ0�<i�;�'>c����ӏ\�-�O1h�џ,����ɒ��Z#�Bl�?XN��c0ø�Vo1Ӯ)�E� Z0����n~($-�?�p���	�4�:�|+p2Ȫ�]�AX��9���Y�X�=���U���æ��o":s+�q����9}<�CB�X����x��Dr�柾�3gv�'O��лJԯ�<m�#b��IS߼e���tI,9�aS�鿶0�.T�{�p%�B,�m��b�����Ӕf�l�>�񜒄�P�d�m�����b3��=L�!cG
���O-"� c
���o�M�Yg��A�va�ͼЬ�78�A+=O&]t%����k��j<_�0j\�&ak�=Ý�`�ݒ
m�'S�a�t[��!���9K���L+A�p���<`1)P����,f���:#]�D'm�r�}Q���be[]�������w�2���I����GA>�P�Q�|�Az�*����3�Ŗ��<�a��e�SG��8��=�����{@�p�VCF+dĿ�����ٻ�� ��v����Q�,.!�_�#]�
�S�/�X�+��Fǚ�*�͂�C�~y�Џ�
-$�o���[��V�r8�8욧�L%+���D'����mrr�Wae��l�ɾn:K XӫEt�e^4c�����wG��:J�;gŁ'g��	�����{�}䓧�w��[mnޒvc�dsw��B�/�M��wMl�EP��d<��s�k�/�~��Q�*Ξ��
�(��Qƹ4x�+ahm�k˴s���?�'���R��L�fzR�U���8^���M�#�fBa�����v����i��9���@�D�l���m��-.��#�:v�����a��7u���6F�/^��=?��b�6���GW��g� �N~춃L�(�Zx5�>\ʣ��ZXÒ8�-�H�)���O��FH3Dr{�1p9���E����E�	y#�?�y��	�"��B[��ϼ�i��E�����=���+y�`p�e��#���y͇>L���X�s�	X���fW-�+z���HD�ċbo�	�c�E.�y"5g� R�TL�7�|��`�=#�u97��H�w�n�_��:>D#%��;�?�޲I�d�:a�q$=��6� )I^�h���Z���=/ N>��>���0���@m�ք-���_�7T�,�mc��V#��{z`ClQ�v���א�GBs�a�=儾��D�)��ϼ�%��k���:l��(�ŏ͊�]}����	�lS#�/�^�ٙ�\�tyAW�c�kINZK7��1��}t!t :?D��-~gm��Z3��4��I�|�9@dp0��vl��o�(�f�N���K,{�Bo�	X��S�?т&���Q�.\�Ը��w��	B$�ߢh���K��q=8��&J㭬����P�����a�K��NT�����y�,Q�<��F��Q�m�L�ocƏIu���x���{����q�wvh�q���(����r>%6�e|�^x�"XtF�F&/A����!�U.bmF񆷺J)O)�C�zݛU��sX��m��J�ص��dNx 
�0=�����\���+8+��x�weO'>�f��*�s᪥:��B+�?���e`�� �3Iѭ�����C�<n�p�KD5p�Tq�'=�v2w�Uaj�ܘ�,�l�t�B��d^�4�s�c�f�nDF6W��tqƋ��V�n��
)h�$7Oub�9�?��SY##�Ν�����*��ϳ@䑍H��G�1)��M��ʆ�ŷM��k�c���F���������v�غ��X���8A0Ryv�\�m 5���;^�ا���=���:��,7�NZ�m�p>ڔ����;ri�Y�24����"��9����y��Sc���m
giP.�^wB����C&�I����gJ�����h&�_Y���߬�u:+�����LǨ^�x��b���,/g� iW<���������AVk���	)c�?a/lzS?D����
�B_f[��
��3^��o�"��
�������%o��A/��$Hf�hF���H��F[,�8�>�ʤ?�
'��;[!���pj�(`�Q�.�� ��>7S[o��M�u51��|_���� �Ę����{����;N�1��z�5�gV����r\�
$#A�<@�,�QHc���H��^S%�[N/�"�Q:;�~��0�>�NtH��a�~�u>���-T2>e_�x�5��8�T�U*��ĝE�;��#�1Q�~�&+���������S��%�P��˓x�Mͤ�r֙��¤p��7�)Q����ث�~H��h1m��c���L�M�Ư^^uU�N���'��A&�b�̹?~�Z5�5l����pa����T�s�0v��h蜭��f��������Hİ��ሁE5�_ 6�)Z����V��=l�	�!vST! 	�k R�!�"�d\d���mN��-~����q��"��x��9���������3���~��g.4�\XL�a3������ti��Ϋ.���j��+�Ǡ��u�`ܶ|ŷM�݂��x(�v�w��$�y�_��m���`xxV0|�¢cE�5B�+���qp
�H���J1�%�ޔvS��n����u�U��s�&p:21�ץw�Σ��1N3��v�[�U,�+���4(�-��b8��q��
�6���	�q�� ��r���V�����z��'z��wkןM����b��� �8��/%m���`v�W��K^�aAĴ}��7�Op�tm��:�_P$�手e��B���K1O��8p��}g�gq=��6�2�p��^��n�k]j�pӮ���q5�X�!��׆`�W��5�����
-XlxVHYEB    f314    1b50�O�9� ��V����o���?T�p��ƪm�s��AR��r%S���������8�����u��pBx����Fǀ竰"��=J*�k<#�j��\�)w�wc7+a%��KG�{�~�PꡤBW C��Ԍ:��޹�&{3��"����ŉ	�י_c��J�0����s�=�R �=�W��dRܬX��������D�]w��xޞ�Ԫ�/�wI�j-$3>��hz�yf6'q~�	�Z�?�D�����Y��|���2���M��k��@�I~"�7{�,�c�ۂ1|�e��yjȕ �qC��D��ܸvų_f��P'r��wu��VS���{I�.[���%^�e������e8.kYه*[�$l����{�����m�1�&7E �˷��'�b>���˩��&:��fUˈ���F���ub��/����6��b���1���_{�袏1l��$��ܣ�w��y{3���h���R�ȗ���~�h����-ܔ��'�(!�&i�!�R!��aE{��n�)f4޽JL��[�G���Ji�>��A4,��:y�	}��A/��%^'u�!C_��ց"oT�N��0��k�R�	�)za���S=ư��2�cv��3�6�Ic#�+Tů��:���I�u^�1���(Y'�"�6��z�0"�i 6`-	��X� �q5�]������!񊦸kT̛@@*0�w='2�Hm��_jܐ8�	 �h4=���GmN�x�(,ٗ.�����γ|)�����y^��`�U�ȱg)~N����4�[�Β�j��5g\%����c�>z�RZ�|ka���I��GoC�du�\,�^��N:c�F������Hpپa��(N�%����hy+��tx��b(_�u�bqo���U:�f8q</r�R�"���&��¾����R��v�_�Z�w����}��&��_d� ��;)4��i^`� ��ZI����?�)�B��h�qV0�G���T�(D���u�`�؂Sw��M��q*�@�UW�i�����pat�%.f k�e�2���(k~`W���ԇI+�HXM5�
�c_�ryoSB��l_��w�8:�Ol���@��1����	$�!Ga���W��M� K�����F�Qʆ^��T���w�0���P����N�ȡ�s�� ��my�zm���@�n�O���rd`0����Q@=�!~��L���|�3�񯳋zA���O�"��g��g����y��r!��q�+A��c;d嵍�j�g�R �1ga �S�s��N�L@/UjJp�����1�!�H*���0+�x��T�~>�J�lRk�I��e�gX�BI�S����\���e�gg�������)uG{�U_�O�+��L��/G?1|,���908I(7�I{J������;#G 4D�,�c~'�1jB��Q�.�j}�lUCD�.��j��ѓ1�,�kS�fxY����H��Տ�(1myMV����W���(?&�V>Ũ�{���`	�:����_}vB���u��{M���I9�,�#��$1ۑ(QG-+f�R.kX7v��Y����L��m�8�b�z�͐{8Q6PT�H��zS��~����?�i�Ѹ�ʆ`�é�*�i"�8{�p����~W�&p0��!mty�ҩ��a�mE�DXi�qA�<�Wrzrt�Nm��u��ER��ǁ�o,�`��۝
��}1�=�UtM�]��FA�[op�I!�e�������u��B��A)]�E��YazE�|%e���M��I�J&<���U�_��}q D�2PU"?v���8�Dʌ��1��1Hm�F���ZD1i�b#'��륧@�"����W���^��".��f�d$�~��D�rZ3k��Ɛ� �ى%���"�B�fT�"�1@�q�(����������y�܁�S��km��T��`G�ĲO�M�Ȁ�C	|�|�����)�W���+9¬oÒ�YC�{J��m��w
c"�*p����P��n���߮�--l_����*�����h�n`�K�Z�	�L������Ҧ6��f\�j����G������>�@�c?7�]A�K�.�@���A�M�U��Q�zX�l$e��b�Oq��@f`JW��^ʣq(Cv"-Χ��ӭ�#�d�ݡ�$ll��^L~����wo5�'�?��{Í�0uٚ����,e�h�����ͅ��81�sX�K�%�Ӎ������&z���Ush�~�k�ٽZ���>'1U%�!�`� <��v
�&��~ޔ�O~�A����xt>+"|�G�%�;�
����h�8��KfƗ8�C�w�%8��:4����'z~�����	����3:��)i��G�´����o�v�ۉQp�����UHV��fwM�ml.Y�\���^��C�,�B�m&<��_���+~>cj�-f��<KJ�w�Dx��TH]f	@�aJcs�'�2ov�A��}�1��/�]/��B�}���s����:��� [�K$�P�^�Eb�0y⛝��K@P��x��Wl���Q����5��Y�V9���}����3kHng�߬��N|��o��ٵ�ify���Rc��ªR�H�c�=+��m97H{w.��^�?�O|to�����[�/�rrSZ��R9��m�A�)���⸌����ۿ!�鵲.�����\��>]��>Y�Y���I2ɮ�ޓGaX��`�����[�>����A �ڄr���_ml��f�&~�����C�ގ�}�3�D��t%�kj�I��6�X���d;L/P�*��Ƅ���{E�٠��Q_����\�� *����)�/H� !sK-���ʠ�;���=tZܧg5܍�+��@4�L��p�mcS@3h��O8L�03]�ݔ���#j/�ڨv��3�����\�����3|A��(��d6�	���E�Fi�d��d�늮��ܼ�{� ���5�P��R!�Z0#G����Rكklb��Sƅw@|����tv�1�iу5�Ⱥ	��>��n]��GN�\�0���>&��h�ebc�5s�J~�{��#����9	z	^�ب>�οZgu���!Z�(��N~���5Gw"��\�� ��!��Q7t>����L&���Ȥ�,����}^B�LH�6/��(kd{�����(����
T�̆"ȗ� �c�W��;�U�i�)y�\oc�z.�<ԫon�}���E�U9̅S;Jn�EPA��&f�<3e��LO[3��?��M*���8�$���,7�y�.~s����+��J�k��f�D-�Ӻ%D���A�҆������˨wa�.�����:��7� �kF�D�N�I5�G}>�~������b��W�r��]��v6-����Y&ְc��cL�,_��p��/��J��0���.���-�]2d�ݠ{$')ÀE�M�:�����S]D�����8��S�������2�>i�:Y�\����	C�X�?*RVv�߱ov�����<*���9A>��a���!ek .J���;25��aJ�dU*�$t0�J� 0R��}ZXDo���v�O��&"�e��������%\V��. ��Y�{ࢡ��Rص��7	Lm��M%mRV`TP#�jh��i@[���ʽ��ۗd"�F�Y����o����_?��쓯Mh#�=�_ه����n?�q��'n��E�|8��mPh��\��j�Z
�*n��g��0Ɍ�uÛZ�45�.Cӌ�ΨN�N�-;#pV�AZ��*|l��]fe���yS>Oo`)� �#���}/]��:�L�I+뒔��ni#,H�Q´FN��z����R�Yf��	X�w���AAZٽ��}RЖ�X�W��$=�>Ip���e:�����@���{cr�e�c��"���<�<8�M��:">a��;��;���_tj_b|Ѯ9� O��8��ش�Wksq�b$�[Ԡ����0`M~���e����J�I H܁.���ח�u��>�d.X��h3^y{�\[��/�d�����g�� b	��� �W �Ї�!A�>�-����O�"6���]4p4�4��Q�� �>��,�VȲ��F|����O����Vg�J�� ��^iϗn9���3�S��m���\��g���~L���۰��myB��4!1*�S]���thCp��s\�>��I.k�<�f�7����~���w�겎D+Qi������q�ڌwB���٩2��H*D�a��C�"���Jt���hN=��(y+��)�cL��GP*�T�a_�����`VQ�@;!3~9��K@�Sݴ��}0�Yt��pM�+�Π�C_S�^��7��@f������?����ZɆ��1c��L�f�k���t�����%Aޟ'�&$�(Ǹ�L�@���p��љ�l��*X�Ny��Z��X��%w���یM��� H��"7�-�����#c���N�����g�)>��.�(�Y�O��^�~�{��V��P��
�<�~I���)Q��ް3�㐣8�[<Ú����n34�W#H�N=9��O6H2��!���n�:�*,�f��ȬȅE�d��W%;c@I<��С?I)�H��s�`Tt��M��}�����%�Z��k�Uc(�籝HL����Q�R���Ӈp�BN!��io0�2�N B7f#�:?���Uu����/�� .��C]V���QK��(~�N) ����� P���O��!*�yߔ�"�"��S�P��~u$8�R&���>8;cή՟�f���À�OE��@R�����LZ z�5tSIpV�t��ȹ�1Pa#P���
�G�!��I��3\�����T���Ѩ҃�VY�Fk�%�/���fj� $
�":���4���PL�����
i�Y�ݚ�DqS���9�� �]gf�QxЉ{ ���wr�_�8�����a������*�2�@58��{AK@����/��nm9*��w��a��=z�y�PǽN�ͳ��vJ��986��lL<��\�성�+ﳍ�s������C��U�8�w��!F�f]93x�]�%��-s����Ҿ�*'�e5�3<��5]�%��VW2�w�v��a�� D��!�G^�w�Z��|O�u�Z�� ��e/,fRy_���'����Wkh%�����B�<Z?�w��g��C��m�]D͇�^�&gq��7�ͺ��D3T�K�Վ���>�H��ￋ� �<x9MKe�0�2����-���dg��B�H�ylzh���R>H,)���d�w�7��6v��o=�!K���Ʃֱ����P��O�㘡�P�ap�����^g9R�vJՍR_��BQ�����-w3���B��� �0���*��O�{��3$-�;$�+}�1CY2��@q\���+b�T �:Q:�U� +y�R챞��LF��%-��v��!?x��+���~��"ە�Q�3;�'|�q�"��Я[Oy��bg�ڦ����,2m��k^�F˭�
��%�In	�j���l�y����Yס�&}�OF��5�S���xI��<�I�]Qt�H�L&�7~ ��?����'H+Y�g�]M\6� 0��'7��?�g=�Eݴ!�&<�T/@�	5Oҹ�2�5�L����Q%��Y��KGZ��ݤ�b�Vc������œ��Rq[�9T�r�G1����*o��m�ۨ����cW'���Z��_]�̺�{~��,���AW�Ŕ+��J �7���z.�o �]��H&��͜n��@�G�38P���aK��×�B�G�(��;Ox��zF�j����'�+2��m�,"@���8�m�����%6.h��BM�w
�r3�D��UB(c�쇤x���8#�}L ՘q���U{���)�z�a��2�x/!�2�<����\i􂕛d����u����P0��-��1����s��� �2k�I�1���b�%�y� ,��U�|Y�X�L]�q��,�\1I���F%�{�B-��A�5��1�9�Q�"+�f����������Y�F9 m`'z4����0�L!`��̋�]���C�T
��}̪,�a�)�[+�v�3�A�;홰R��$��oF) J�`�p�Fj��Mp�W����pt|�@
��Za�C��1����Iƫ|tSF/��W��J��S�ga���0����f��s�#��N���C���	�%�ѣ�5�����X�G9�����`P����Z��8:Pr>DiZ�E���7��G�lG/���p�u(!��U�ן�ì���:g'a`x9����С�k-0Y�D1KT�&�K�H#&�� z���.��U�&�`gTJ��l�M#WN�n���=��T��JtYU�!\���V]�oo
����Ezi{y 'T���?܍����x��`�Q��To���q���Ob���=O2	�;����U���t��#�R!i�Zr""i2d�>S`xq&���^Mj(�v�g�,pem8Ѓ�z���+�
�� 9H=؝y�86JR-E��,�>S��a�KU.f��e�˞e���'1z�k�8��@������_B�e��[|0-��;e����Y~R�O�w�mf����qs^�j��{@O���G$4���u�J<R?�M 8�jO�{n�x�"��I��_�3�?v������o}� 3ZAs���dӭi�vŨ�mq̪�1u�b�"qv�(���!'I~X�!�j�}p�U%�ɮ�D/��H8}`�-RSǩҸ�|� �jL���C�h�<���8��&��8\퓄r������#�g����;>���;�m����� �.�ڐ���r�<n=N�U��@�ؓ���`k��Sр�7�fF� ���[
��9'H�2��f���C��G�Uq�>KDo[�c����s�<Z�