XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3� e�j�5�/�,&���b��F��t�jR�X���\��7Cn�����~�q��P��R M�#� �:6��nS�ke�j���3].�y-�hf�o1	���!4����vG�:ѰraO�r˜5l�_��Hy1��[#f)���[8��t:��+nt�.���C��G��Hr~�c�����?�F�|E�\�m].��쾒)�*w\�9], �L�gX$D���h4���W�����~d;� �p�����R����Im�\�fŤG�L�>�0C�FD��N}���"�r���Hu�$�����A�J`JnK��߫��t�O2aˌ <�2��{�\��E[�A!J)�t�{��Ut��l��A��S%�͋L��i����>����#�#��
�+�zA&��J�_i��2��ޥOm8��k��C��P��y!V��f-�nj���
Y�<"��S~�{X�c�	�{4�;b6Q����FY��[��x��K0�K�A�:�T���x��m�t<<G�'̬j�;p5�;��M���� �����_����u��Cr9��ƕ�U�{�+V���z2�֧y�q���b�v&XL2P��������+�00��e�����@mgX�~�s�F�>@H��TP�!�i�Q�P����, ���|.n8&��w"��wiΗ���t�v�Ÿ����m05����O����K���>���G�t����;+���)W)�OC��NnײΜge |�XlxVHYEB    fa00    2030g]a��Aʴ�Bfla�N_�E;g3c�5�9�����.Ͳ�m�ٓ1���ǘ<���8U����Z��a����9����/�,:i]t^�W�Og�ޘC���
<K������}���K��	m�M7�Y�S���h&��	�B������#��>����a�o%OF��,5x����]J}L�9�t�����9���-[�?#B��xߓ�1���%�6vj:A�f�iN�� �2j�S5h���7W����|�B͕��8�&�ױ��[:���v�'5<\6rߊ�W�Ҏ�:?��}��آ�G���zrWtn5s���-k��s=��t�Y�q��O��z���]�맷u�4d��K�U�&_���l��-f��3�{��A��r��ٔp}�9i�d�#���o`J����{��$��{a�Գ� |�ȍǓ�=�Ӫ#<��Z�h�q:�,G��q�L���1�*,�o&<s<���0�p@=~���E��w&�������zǴR��Ї�W�N���?�gS�w�-fR�vI���$j��g�P���;q�Q?g��6
��<��4�&��� ���d��E\1;Đ��x<���@�Ή�d^���(��:c�V<�d�@ß<V�BbK�&g��S�ۻ:��[�V8<��9�\��}���&'�����T��OǕ���R��-�|�5�x-1��9p��r�6:C�@H�Y��^�h��e�2�e]}Ҿ�d��$޷+b6p˞~�h�u���n�8���k`�Úq��m��Y��v�;��Y�vg�Rpaf�7'�e><4��6�t���;'2$?���~���zy�-F>�y��$�Y#-�1GcA��W�H<ջmQͨ�$=-�_�	�����xc>
���>X6"`5 �#"@A�����)F=h��G�tX�3v��:�$4������R�:����>ë�`:�\V�9XF��2��T�Qp:O!g뜿.QЯz�Y� �x�X��������OW�y�5��t���EψLA7W��)�� &c}����L�Q�S#��]�Ӏ8b�N�+{��k.�xl���d 
�Y��Í9���wV&����7St� ��o��\AR���?*D�����`�慛=9NϏc���K��� �20�������uL��X�e:c��̹U��Y%Q���$k�ӓ��D�E�z�>mj� ��<sR���Y��y���y���4�M��IǗ38���� ���?^?5�'��{�՝	���V����~=��C������fW���A�?Ќ\˞��1���o�`7����$�����h��(��,���$�χ�v�±�+-V��W�������2<uץsI�R@N�*t��|'��-����R�܀���U�ٷD~-#q,������}������,����0���C�3�R�lE�<���X���g�9�M>�� S��Q�S�M�|(d�΀I�C�:�Q>���ӛL���L{~ӮU)�
 prk���(��Ġ2����wA�A��ď�+��3i[�ѓ�Q~����Ӳ�I/���JK��L���^�ZɁ0�v1���v�5��I�u���gi��z͗e��\�@��O����_�<�;K[���X3�J��_�:�^���=��ʈ��T�>l݉Җ𷙨v�NO�YhcԽv��$B�s��q m	��;��~����V��Ɲ�C����Q�	c�j&M�.s��1W#V\	3=k��o!p�K�΅>1S�sO_t��n;�f�J�&���lĎ�������u$�D����ˎDƁErkL��[o��<�E����P�U��� O[g�6Wz���ݘa����k)�n!0����CJr��x0�FMjw>˛qUF�ҭt\r�K�e�h��6����v�+�pN�p��d�#q�*��X���1"K�|�~�#�.r�Ø���w��a[�fh��~�b���%�K��%Dp����~*Ӓ�A) 7�6��ݨ  ��j1����͂��X�P�>i#�$؈G����Ga�$N���ȼ�Xü~����ֵ�k��쌁p\B��+U�P��6��6"f8O�SY�*�����z�4il�>vs-B�g��E�{�ڕ�*�� r0�hC:4o����QC��s��m�+��~4H6s�Mz�n��J0�8ݓ@���<��^�0ҥ�ѕk/}��֎�o݅�8�]@���]Ha���-d����_<!�96����@�[S��lI����'�Tϗ�����86�|��N�7�=*�G�'wӛ����9獿��b�sO�g���Y�7<Q�E�NL���H�_'�Xon[�����3�Ř��A�)���>�*�77?��M蘳�",�G.��v��?�����K���!������ip�v��Pּ��D����gT#�hUw�HJ#*ۣ@H+An��%Q��a�z�����}���J‑�R�Q�b5�?&ӣ��������F�1�Ϋ�H�Y\p�:w���*`���V��ﰂ���
�,���v�b�&�W�
�ψs�]������d�w���fy�\<�k�8>fv^{�]���l~L_��R�Y�$����H۟��u��٪�jk�Uoj�ېIG�~�+V����|�*���o�^5�`�ٸ��M{C7�ϸ�h�����t�6���5n�.���hE��X"��U�ˣC�ѷ�������m{b�ˋ@�h�#E��?�L>Du�~_2��8��u����C>Hy��8$��-.�|�k�!���.�g�9Ƀ.v;C#�Z�d��R��X��#��\��/�����$���api�)d�2N�ϓogX�k�I$���\�����i􀰧��6��栤�>�(��6]�����]�?�uP�r�������Y?Iis�m~�,��v_�N���LU�8���� ,U�J�{(��r�|\�?Q��F���5����%֜�r�p��CS+3�i�uf�O,<A��|1١���F�?�d���x��.)|V�.W��>�V�k�Fb�v�N���M �G�'u���*�c6׽����B~�hQ�P�[@�X��mZ/|���?��p�+G��M��W�<�r~́0�(�u�8Uċ���`���?ހ��?��w�57�#�ϴ�b�]�Y^k���K�w�µ0?��&䏌�4>��f#�1"�d�ˢ��r�����A��ͱ���e�!x�ݹ����hv�w|Fɢ�<�~ї�v&��(w˲R#B�C�r-@�����f�~�0��y��׷B\뙸�*�uk�������8�H*���o�fr�fe��(���~��tqE�����n
޻>��7�FP����s�[��X���U���g�~���(�i.&�=Ɠ#6eӳp��ĈEl@6Ѿ�'��3�Tc��c�)R
5ߡ6%�A����e�k^o�nؒ�#x�VM��-�L�\32��T�O����[oz{3�2F�o��?p&R$�G���Zx��\��u���P��Zk����ȼ8_��1}ؐ����c��ʜ��1D�. �dA(�XD��Iґ�SK���9�YGR��(�E����iF<�Ms k��J2���F~1��[��8��%CN�o�S�p���2�P�NhFN�����zeP~eyYL����LO�&m�4�v��0㱌��5U)�����d����N�MW
ڊ9��G_xv�:��o��'��;��f�S�f�yi�,��s}��r5���������L�"�qt|���]�Qf��5���;R[F2	/Zu�2� ���%�L��Գb��^+2ᝈ���;�|;�'��=��RG�r�7�~��=�������36&>.';쀋�)�sFsp�yt��7�/X:�/Ꞽ̧�,C^�(���~Ca��qO4��6v�&�����Wc�j>j���3�[vl��z�W��>�%zĮ�UOB+��M8� �i� �%vE���ںG���z�����k�����|�,�><#��~/~I������@L����#DM*p򰢶ch���/�t��!V�����I�ʿ�yh��1�^[X�¦���g�uoJ�O�(�����=Gr��H�E��%�6��Ƃ)q���g)�PldmpO��d�x��K�p� �-c ь����{��ۇ�T�u�u{���-�A�	+}~������w�d���](�o	/�wѧ��(�� $��cN���S��Qh���Pb`G��6������ �36�rz�-�д��bB-�qh#�kQ��qO��V�;�꘯�dI	�[AF;��%�mg]�b�l�`xM�_��I)��{�2ә�%smrV��
@.��-o�"�%z|�}���r2���d�=�]�
�vB�-8�ޕ��w��R���1E&�ȿ�w�ٟw���OD�г�)[��Ȏ���4'F�\�9��u>�4$��W��,�$a\K�����9��^�v�}Y����y
L�Ht�'g��d�ql)(��N��y���8����j�����#¾�2e������{6�☙z�e�I��r��J��;:Le��9:nx�m�T37'����거���p10kJ�^�8`(�O�׿�L�8��SK.��V 
s��O��|�؄���5\�؈ކQ�	t�c�{o2�K������"˸@��l�]r�L�3���6��yӦ���]Z��u[�u�|���P����_V�U*Cp�y%G$N�@wU(����U�O�-LvQ�;�"��ϼe^��<� щњ
�2�1D��誛׬�)G6���H�&�@�``Ѹw����]zCW��'	�X58F�?0&�_^yѿ�闝��N�{*
Z�8���{&�5� 
`�rf��8�B���M�~���Fqz�����N5=��4_iŇ��3Vg�V
��X�O$|���<�=�^���c�e$>���Y`�Q��^":����z�l����UӬؕ�љm���b2�.�@�=����}T���m9���6a���!���1e�a�s~�柄̾�"��n�=qT��ѫ��p�k�%�)h2F�!���i�5m����ܲI�BP��HP�B��P4�U��%�ĸ������FR8�HN�v�j]��&�4�	N'��� �o��jWH��H��RP���^����~vQ�� *=QO�Fh0X�߹c��:���7���� (��|+4RW�hv�������Qy�95U``M:�Y9����_�|�#M��d�u���*.<�c"��VC��O���{�O��pl1�p]��'�K�EQUw��Ё9����3�c���P��z��bh%�� <��<�G\���q�æ���3V"3��	��ن P՛}������}v]��30���:7�1�af����'G+qy}�
h��T�H�"�����V�愴�:C����K�My����z�[7G?;Og��`�'�(;��o�;B�������U=�EW���Yfm`<J"��Fۙ�L#>H���T�.:W��4a.�N%5�#�DS�N����Ю��K���S�/)�2�y�R[o�.	,s��S��	;>��'�y!t�k���f�o�^�����W��/Z|�+�1M,t���V��ޛǗ�~^D��-`iԌ��0$ta� �caX$F���8o���lt y��a�ٲ,�y��U��ѩ7�H_"_U?q"�m#]�n�s(z����7Rb%��Gm��������b>���p.-s��#��M���8L[֊w�v��;ʒ��ҌJ��tjR��(�	^r��ﶓ�y� ��� ��:ݎ�Ԗ�p@�6_�p���6o���$5�#a:q*ʇ��3)�O��Q��A�~�Ex�\:��s���vE��ށ�h����"
;#o�F����!2�g ���>�w�`�:�:�z?)�[N:���7�'����HeO��H	&g�Ӄ"��W�!��D����?�<��M���ҟ=`��1��R>-�	��_��)�Y���{��8>�D56�GIn�~'߲���h4��v?E��u�nW�'+|ōˊ���<'���"��J����G(����\�G��S>��㸫�Q{j�X�a��kp0٧Duk�#�ʳ�H���ؿ�T������v���3���'rԦ���Yt��9�P�-��׷$p�9Kwz`^��BW �-'9��F -�`��-�?"/,�;�8�6#ufu�8KQ�m�L>�2n�l��L;��bLT��,��!79�zf}%d���C�- �xL{_�\Ѽy������yg�Gxt�|7���$�)!��?��R��ܑeYf���T�78d�]���׎�C�P� ?[�^Y��`�:#�'L޻��Q4hm<�6Ѵ�c���5�c6��m �%���=A�7>oI�҄�	�e��a�m��L^��~i��1��e�̫&�㗒�B~��y�3���ʱ�Q���U���kuk;K�p���|�;�O�[F�[A""����J�$���z��j����g*8i|�Ъ��<8I�F���\������?�|�h�3�n���K��qЃwt��5&�h�6�U�JX)���aĽ�'n�_�|TE�I3�v�.�f�\]km�]�b��V9A�MFW1���`�)��ǀY4W(�v�$��%u!�WՐ;�*��RF�ݭ����JU??�;�|��-�{8�/���o�I� ���πS��L�=]'���!}�*�����D1�*o)�A�Ȱݼ�����d^V�B��!��3�S6}�(3�L�9x���n.j��r�����xn�FN���F>>��#|4<�e9��/�����Yy�#��;I��A�:0]a~�kw2���8����)�r����`��q�tr�A
@~�.�#"d�����s�+�̴Ȫ�9��ʡ��MM�a��4Լ�&��G.�#	�6��ƌ�O/�bnb�Yj���GOgH�N�����X_�Sf�qJ��~~l��z1}V�f �>)d�~����'Ր�KN���+�6+��&@T:eDvh���������,�(;�P:���2�����n�] #ךק�aO����E��.S���瀻[VU	��п�]�������S7K�\Շ�KL���)U▇�LC/\��VCjy���}�te�Rj��H{�.v�E��X�Nm�T.w滄�a��c	��8*�aE��ޓ�A&Y�;M�4���sy#9�n�m-�[�}'9�`*�V��≃���9/E�&������T�f��T�����o�s*�)H{��*����8;\j�R��6�\�vWR���	�U��ɾY�a/��Ջ8����+��1ݪC�O�~aε��]�aQ�R��S8.�xek�Xoh�(t�S�5��"�L�[��v�ӛ<yZ0�/I�9���Ψ^���tQ���'Gz�G)�As�Ty�7�뗪BN�_٢ՔX���9ʝ��,�|�B.]���p�f��%Q�rZ��_���e�g�!��z	+���e����U��D�7	j�����#MU�몔�>��D�'.�JF��K;�����`�<N&D��6r���M�Ī(B�ܣO�s�����7X���s9l,��u�Li-{A�nQ���ߝm��|cq�1l]	?�7����t��±�����O\���P��x��@@��b���B$+X��{��A���c������B����fΥ�A�����8��~k�6�`l� �6pi?,��ҵ��Z�7��+��o���t_t�SI�-�*�������ۛ$��'�g�;�۔�K��.� =�c��K)��缂�:���M<E��|6�urf�AOD�c�$�e�[����5X#�{|��
�A�{�ԛU��0������SZ-]M�R���q�5�*��w)M#7^1-?�s�������~��	�^�5�k�Zx��Ȩ�ɑ����n����H�o��P)|�>�8{�w��]��/�b��G�����t�I��L�1�0nE��~p���HKWe[Mǐ�@!���;�I�(����T���Ǘ�m��ïs��e��o�F��f�QU�jd3�t���%[��ϔƾ����'4�Z�x���K\��mfD"~~����71P�����t��8����E�+'�~�d7�S�*XlxVHYEB    9620     d70�a�m�
�$DY���ԛJ]I����)��f�#����H��& nM��h��]E��Y�_�҉���*C"��z�����8�]��1�ĦP��moj]cN?`��<P��YGh�E��=W�������~�����$�꫗��,�K�I��c��3����>�y�"���n�V]�[�nV�vX��>��ZW0?���z\��*�N��
�˚�P�"�B"p�0�^�f�/
��<v>���ቌ�(h�rTG��( xY�#���oC���cU�&OW�h@��d����hl7�������|ĉ�.�p�S���
^9'q0��<q�H���?~�h��'VH��u�/�c��N�����Z4VI�U�� �$co�Oޑ��y�d{��"П4�h�I}K�괒���(ւ�N��l��2u�ߨ�#V����C��DG\���G'�W����X����]���-t�Y�qA��c��J�D�71�׳^��V3Ҍ���ĩ��|����� y$REo؇c���!�:l��@7��L����#�|�h��o^�YIF�F�	���53$�k�xʙ�>����^~r�赜pZ{��=Q4�(-b8X��<� l�α��yO"�z�I��b�;]��R�1�g	~��-�FuYsWOchs2hf*�]��R\�uZ����$wq�!�n��J������a_���2��h?)ݟ>�p�sK���E�g�AЙ.\������$,��*�؁GZ����WQ�r��ˤf��0��VŅ�r��xt�,3R��-{M^�7�$�Q�����d�庒�N�{�����w�2�0����j�����Ny����s�V��k"�l�����>�pqq��pf����G�>p3�Xw�Yfg���E]�y��*��ɣuw8}Q�CJ�"�_�.s�ف���jA�u��G{:䈜ѧ�_`���4�!;��H����}�;B\��Q�QAH���E/ޝ>�{$7-��ާ"�C�ղ��y��^�s�4��O�Fq�%��S<yw�G��_����?)5�ґb��D�n5�JN �PKJ�-�p����1��/ߔX�v���:���J���1WlI��D�����4��v�U����?K�k,O#6���'Z�|��ڬ���¦)ST���7,���UXi�t_�8.I�d��H���� *���S����~��^�|����]�b��`@5�1�PJؕ��.�/?�,�b��]���I����W1�@Sm���d������ ��tT��K4� �=�k������N^|: �0?�����_*�}@�a�6��N�J�!D��j+�
�"����v��a�T�K?ٟ�'��VGCE��+���D�'�u�|8+��4a�b�\h�ƵD٫���9P:8�h�LC����v�5�TS�t��$�?,�pZ��xyzR�� �?`+��y��<��Tg=B\����K�8�5�MwH��:�MP����B���D�ޔLآ�J_����@�����1q#O-��^w��3ҜO�w'��]�"r��<u�j.�K������q�ȍE6:X�=�إ8�y�@,i�G�?,>�t������ҋ��\��bkeL�(.w�Gm���s/�C�|����D���n���9��-ƈ`Ov ���E����?(���G; 6����U��e��إ��_�ĸ���¼���@��3�~��q��=cf߽�䜁ɴ鼶���|�K��'�
�9�썄`�6��H������=��7F����z�"�vl���\X��З�3�o`lV��i����S�9�ǟp�(��y���"�H��k�r���N;�/�ЉX(d�D���p�گ�J�����DH)~/Ϯ�:O����	�0���^@dI�{o�f֮^B��8�;���� IH8��v�i�/���Aםϼ�a��\��h��}����ó��5�R�Y��g�]4E�`�O���c�����:A�=pT��k�?�IC���hyw�%��ʀ�a��齊<ft>�_R�V�\XK}Qz�`����)zb��UJg����e��TM��h�f�����uB~=��_/����J(w��̞.#E	iw�~k|kE��ˀ�$r�������Fa@J����m�BI��v_F�Lz����(@7
���~���D#�c�W�ư�Z=v�@�[Y���ԕ��� �������������<Pr����� ��䫭{R)�{z=�FL�s�1@�LCs���^h�%��*�o!�������WW���נy2��M�׹��,����1��y��~���G!	���HR�$N�ˣ�Ί��uO���~ǍRﴣ<R��J ��}�?���~H3 ׂ0\�س�4�[�f��%���ꥒ<�g K��j�Z���5���#���,#���'�q�6��H�����b��󀅓�����DT���q�D��eK�G���d�#s7�F�t� ��p�kp�B \��Hj��s��i���w�f�\.�D��.�n��cA}7 �N)��AY���b#�*��+�r�ü�_?P�ĻR�g=Qağ�	�<��i�9Nxˇ�nd��ہÏ��ԧ=���|�?	��������c��4	�"����l��v9��Lr���qU�札?�6P �!��F�u�~���@�\N��S�i�p������2�_�0�Id�!��<����(��K+FR�$[��,���P��^:�D���<�7�����pz��n�-����9u�u�i�j�Rs��L��aL��>�(�
��*o]�e���P���X�p����k�P��,x�I��ʤ�S�]PX
*�Sx�^�t۱����>GXT@�t�G�Q��%��t7��Mn���qq����,%����Uǐ)X��Ԋ�;��v���L@����S�GT?���н�n�Z����	�v#�4�S{D�����{Pb�xp�Zs$�v[��{�x��w���jF��U�V���_@AlʨVJ��T�ѵX�'AY��HA�b�0??��ǯwF�21\��39�벨���󙩣-�E�PF*X��dP�N�����RT^v81�[f�);� �V�|t�ˤ5�[��hT~FQJ��`�޽6�<��	lk�.�ETƺ�"�fg�~��twGh�Wp�ݦ�I8�d��(��%a�aB�������t��$�K�'V�9pGE��/i7��4C�p�h�v���.��fe�x�K���Yh	7DN�C�Ry�mI��q+��"Ose��Cg�!�mM0�X�+)�?]B�^���D@����a��2v�J�1� ���}����Um��kvE�#<n�������^Js���ZC�}�	l/8'��!�e��Hré���!�E7zF�+�/x�f\WD�<H�/�-"'�