XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���z�K}V�����;�φ��[03gL�x�>�_c��t�[��
���y�5?��I���^=��'�����.�&��C���@AQ�s���L��4!'5�� ���8���˿}��+/ʔ��$���j[�6���E��4��������[����>����v�J,�N\��F��w~�Q�l���I9�}��6�y��م��w�o?���`�l'j� ���88���jo+sS�B:7�T����'�}L��!���<Z-�r+������S�+�~[�3����#·wu`U}��u�^3I�!�X�$�`$T�r~^19�,���9XgQQ��ٞ�2�%�u������7���B��U��d����0W��X��:tJ���*7�n!:��%���e8z/���=�j4��䅱��P#6xsF�U�-����tI��p7��_`nIf뚫2f��L�zA�T��v�F�~�9z�_��z�[�bO��.x���nk�i0,B����@K�������&��zu����i36z�[��ۧ4#2Z��">��ȱc��R��{���0���8�e�o\�X��m�o�&�K�C�Q��z��,61]�yF:��wu'�ۃ�C�"x��
A�z4����#40�$���͎?)"2egl0#��y��kjX�7P�F�m�Rw�R�!�/��n/-�.�w:"x@�66@�0(�B�[��ф��i��z0�.����ɧ7`��}��(�/e����{�O��XlxVHYEB    b8a6    1ac0R��-�_{g.򪪇�c<�)��f� �B���x bgp�
i�=�Ḵ����Ŀ��%�}�;��|��+g�'�l��6��9�Ţ�K�zx����i]C�R���]�8~�P�_>K+4��|�2�� �x��Z�`�h�����;�����z�O�</��2�Gk�c˓O��oct���/�Xh2y��#� @�y��p��9��|�Av	�g�)��6,���,w����+�R��\t`M�2.���YV�l^p��˙��G������T�3V�A0o������O���h���l`�6��_�AR�[�ͮ�����g�q6F��̳2m?�~f��u�ϕU��8�?�O��p�pXoD��ʑ?i��5T�� 7d[6)T�0�EdVv�#a�`y�,�=˫�����;��F� i ��F����s��*���w�sRgZ�֧�Kn���G8އ{n��_��K�����E:����$nnt�CZ���9�㬡Q(:�j�n�� B�xų4�HC[��R�Yf<Fb)�1���K�UD��JB��=�bu%@^jn��LR�I*�*��GH��{�W���8\Q��t~&�􎔓�E�F�7)@���c���ܳ�(ɪ
cS�崫��Pa�z��D馯Ao��_�)"T�r;���()$8$P��c��kT��f��ɉh��%���Q
5r8����c�L�JN��r{��	9�`�x����P۝��_�����[�k|9e��8��M��^�����m��c˜Ŝ���
��~)��z\[��Ӝ+�J~Ҩ�y��^
�为|y��!��GC�wO.��o>ũCS^�蕹�	E�}�rYޞ�s�=���0�$I'�-ua`�t���ӝE��/d8"��M��I���!;s�S�A�6�P�o��jD�f�f�gY��]��S<�
4Y����\R����8j��(>D��
MZ��߬D'��ၿ���0���ՕL��_�<>C�P�'3���S��D��6�;7�����n-t�v7��EP�,���:� J��u�}�Mːܥ����uWʲ��!P!������5�Ģ����鐛��~�7�q�Z�xG�s�2ye� #QVȘC�R�=��������E�t��A�"��M��E���v�:�ÿo7�J`P�,t4����{mk\K��T�=�&�g4�&���/[�w�EU�_�H���Vl>���'wj�a�"������a�r4�j2����[7+�2��f��*!1�P_H�l��P�kh=XG
$ú)��A���5�*7�*��}2��ˋʅ���z#�>SW}NѥJQ��q~{�w�˱J�r9,���"m|OgDҮ��X�@����$U4]b��L9P2�pB��M�.9|�����p^|}�j����lq�R��Q'�%.=�|�W�^s�ԩ�g��q�³	9���Pb,�l5��=�s��95H��Ȝ�p�B9*	��I.�^�FK�%����p(�e�r��-F�w���e|R��H�B�v�̡kg�����Ny����*� �fc��U��D|����ҥ�G���jo�*`z�z�۵q2����nw�W��a��L`��l�lʈ��o��~(c���S��#����@�ЖG[#v�����b�U�$����?��s���>+ޑ����Z�!1{��0������3�*����e�{K{�#���@8�̱�!��@�S5��5��PnD�pu�C]o��0߈@��k��cV�zO�ѝA���GΡ�n�y��!C�b�D�н�bYs_³�j6�\?��^k��1���9�.d�w�@ь�5�B�� �����r�����j�O��o�������n�����5\�a�J����`�&�昴�C��s�g���t�MJޫ�%Ag�x��?�7BgCw��Ր�s��Pm� J���f� �gR����a��T��Ɩ8��p2��8�W>QLQ��k+��'S��S1~�4�����>5-� �L{/���l�J��F!*�G��^���[�7X�㴨�4V/=ꌿh�@&5����m'ܵ�Eb� �iR"Y��J�MmM����p&��֍n�W�K��0�Y�V�l������5��S�t���E���<��ڴ ��a�� �fҐ��kK���A��-8"�!�y�����CY{wj�6F7�-a�|�x�Q���r����Hňd���F0�Y�qx��M�9�ɇ~��/~��Z����}���%���_�
7�ށ\Y�{i����)�D����89�21�Un��rm7KE�x�s���ǿ�%���s��:��uC�l��҈�P�<Z�Q�yQj�^A/��"�I{<�_ū#�u��w��t�/��&���"`0�eW0�dP��Ƴ��(�d�8O0U��M_���R�=<-{�I���	A?!Ͷ�w��!4����S#�\�(��<��@K:pѣ:=[�>��C��W�͈������р��3g�iR��A	���~宠 ����U�3�(Fh"��e���&J)ߪ����q��M�.����j�f(dR@���?�A����gEgC��f� T�(��4�3l��X1�Cl����m��״�"������S� &�̐�3��ǀ���������=|;��#�H���*��Q��	9G6%�����6���mN0�ٮ F�w�[��ՠ6,�*��ha���r��y�k8����Ƚ������j��`�����;��>�}�Al��:ͦ�D
ʌ��b�8u��¥3N�t�*<�� BU�b�4;���l�z]߉ݫ�|�Cs/����"��]^�L���~��zA�C��:���l�ǫz;͙�W:��Y?P�@�~o�^t�
n�o%+��ak��l��iz����O�M�~}�b���U[W���o���Լo��5t�a��ppS֩���J�J�~�=���W!P��;Z���(B���A�>������Y�ho�J�׋٢�tW��|Σ�;�+��W<����&3a-A�^�m��6���^���}��UB6�pS����p>C�����4��2u �C�dMBQޗ#!����7��%u��ַ'�o!MBF�?��PW8�o��^K�&�ث�-oHI��n���xz��ɣf�q&
�,�P�N/�����'�7��BK����]v�wj�8 ��9��#�oT�
���a.p�[�5������z�|���%i�9V�zJ����?h�6�9��&y5�#�g�u0�[
: b��z��ԁ������[������5���l���7�@'T��F�#��� �%�����mDޕJ���X���9��+Z�!L�.Lg���[�ڢ�U� ��t�R�bT���B�[޹Q:��d��i���B����*������V�o�X@ڊB����&�9F�+���}����L��6׽�Y\;�aYk����勔&�[o[��{��DQḊ-��!S)$�=�h�[�?�N�خr!��[��CMT�Iv�E����N���'��f����m��*�a���h_3#�k\Z�ΙL����������x;P|Z>��!|����q�4{�˶�����b�~��t��>���l���Y��s���G=����<�5p�x\�-��Q���D�Qa#�|ml�# �<c�)�`_H��o$������n�w佋&�j�7uW����K���f8V
y�2jq{�����ొ��uKX�'�֗�Y�b�?�6Y��l�I7��g�`)��r�*�_�#/����B�W4⢗���p�/wY|��S\~��4��d��H;I��1,����eY��S���`z���#e�;~!��P��f9��K��+�EH�vR*&�[~���=��(��M�/�#�����d2�蒓T�����GyW����^�%:6z���h���9���U��x!Shx�@��T9uK�sv	V[I1�q�^}���b����GW�8>��sL��Dy�����`D_:S0C�+T]WB�WT�|��c�o<[o�\+����`z�Q k9���w�o��͜P�_(�\ٱdNZ���{����%���5�LE){��h�l����WR�ȟ��R.F�4S��|>�D�-���L��H����|��I������n-� ��Б��.�;:^WZ�5��g�O��l�%ǼyH�
K����2�P$����ǭ��.e�	`��|���z9�e���*Э$.(T�	�/8��z���3{l����V�p"�ڻD��[v���9�E.�mp�����'��;\zn�fae��hN�J̏+{P�x�Tv�&��S>��!O�0�<B#�/��-j���φ���c���&�,S��F�C2@ע�gDݜL�J�mZ��|���6�) �N�n÷�9gf�+6�?":6l�7�DGEK����v��ML���%�QC��>B��'$@�%E,2/�2��M���'��V;,9�;�H�¹�]X��s�g|�Ԍ
d����/�'zC9�T\�*i�b�W�Y*A��r߹ma!��%�>c۬���N����"rm1��;ͽ��27LA�eO�@L�N`]&|o���1H�@��U ��Ǜ��9��k(d��:yO�y[��b:�_7%9{��a��d-S2��E}�ףN
�|�#��#."s�PX���֭���_����s-�L#�o�1<�Q��������:�E���J�\{T'o�HE�Hơ�֐F�e��#�u�r��0�8��F
�˴���M��x�8��v�ba�Ĩ]�#����\���=ߪ��a����6�aޖ������'0��]9�w�&�3��K���д���90�̀��ӅA�AGS�^}F�|G�%�!c	��:_�aXs$����fR����/)�cӨ��+�0�e�E�X�r��w�ӈ̦X��U���̩7��
j"6�
?N\O[7;-̑�|�;���^�E������b�Z������m�wϡ���+�q8T����1��5$���H[�J�x_�-<E��n<`f8p!�8Q�}N#�.��ka�Q��gd�G�4�P�@j%�JCJ��J`�)'������$�Ut��9��S��$eEC���I۴ �\A7X�ݏgz/чߛi������y�N]���1��c��Fb,�u�}� ALګ��	,��m� �3�c��s��+�2<�pq��Ѥ^�{�Tۺj؋x�i@[�	.J�V����p`E%�fh��Ɲ��z�& 6�rl���}��7(V����=u�s<Zw�\D�T��a��-�I�b�Q�mTp=���_e�3��~t��>CG<�9x�/���5F�^X�E��Ɋ��ը���fx�V��)��]q�D0ec;��H�����?a�1�	L\�-������M��DP���R�X�{��f�V�`��㠥P?^txJ�@���>�B%S�/�k�?�����2��U-ɠ,�X�4(����Lv� +��W������6.C�ƛ=����B�_d�b�Q�e,��0z3��%r��z���R}5DD�dQ2ݨ.U����3.�HRy�+)������C�@�GE��{6�|��щ�'����D)={�c�;"�-�`�t>�7�R�̼_0l)YqUѶ�̤����z��=>el�P�[��u��",
�r��:��>�W��4�ܿC��+�m��(4�(+�\J���UfH��@�g�ِF�Y��5���ynN��_A΀���X���KT���:)��&�XՎ\��ӾZ^ao(U����K���:mq2���.�<�C�� R��'�]U�ְ��{^{�5]>z"I��׷��,����z���05�9���	�]�g��;�M2���޸����~2�^��TB����GJ:�`P�E�S��"V{o�W�!p6��`�:����&8₻�� �����L�I�Ș����	͖�v���Fy-�!�1{����+6�;��/R��u���	=��������`K��	+�� %$�Wr'�e�!�LBm�^�e���ά��]������Ê�{�-=,u�>*%�S��t����³՞i�-���|��11�G	D7�t������B���ᕘ+>��{V����%�t)��u����0_-[� ����[�]���̗'�j&l ��f��I��`{4/� ��g�Q���&��	S��Z�lP"Es�Ǔ�#X��B`��=��TI|x�����k�}`,�&�~�A�t
 �6��6�Oʏ�l $�')M���]�{ƫ�J�TC���D-������s�+��>���[��Fs�2�y-5�j�}MM����0ƺ���G���źv�Z&i�}X#S�w�!&��	�5o-M3�mh���� �ge�0��k�0e�LN}����/KE�dMâ�(����K�ܙη��� _ҽ�qr�[Qٚ�!��O��)(,s���=[;����.�V�f^��dSyÞ+Ml�m��4\�S$
��o�f����͗���>d��3D�q��L�e�q'l�6+:���$*�Y~
dL[��UKψ�C�g�vO�P\ ��sǦR ,k\!�tO���2�C��P�Ȱ������-=��e?_�Xa�n<�T��rɧފRl�c	"��FGV����<U�ґ�����vm�!���L/�c�?l�]-4��)/��N�m+KҪK���ٟ_�R���G�Μ���<�[��߿�y����Q����ы��ӱ