XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���4X<ȭk;y���O�TE坓����&}B�*b�H�]l-2���ȉ�P��������T\��
B�ډ�1�9e��P*�tw��;�x���M�=я#���z�v
��G� �����E�e����%@�D�s��Ԃ�M��X��T@��n�m�g����r�L�ϴk6��FM��c3� ��b���{R7>���� ͒�퀤���y[�ߥ�B�ۯI+����V�u�zR��?��|Xs;��W�g&��o{��"R��r�@��4��f5W���ю��B�|i��+�*#�bv����P8N.�1{��3�"K���_Y���}��AՊ���ŵ�d
A�X��;�I�X4D�J1(��Q���C��cA�O~v�B?/�� u��,�>j�	�#��%8���gFj%2FnR x2�n�bY�Nt�\���V�X��)P���;	Qj�a�Z�ء�a�"��{�<"ѵk�8	,�� �?+Ӳ%�Jg����;:o����A;u̡o�4| �:NUC�EKH��غ�U/e��O7V
�n�8=<���I^6�.� �p �m��� K�6���~�V��ғ�H J}|�]�4l�:Hil�6��o�&�2�o�p�	�9hw�Vl��h(=Z��]���c��3�T斒��۾��]�#<�
�UOM�����ĺ(	�ı9s�.�24_�Zu����T^��K�ƙRL!�3�S�n+�?�	��ܶ��m��$�8=%q5~���ܧ�!�?����}������XlxVHYEB    fa00    2480�w˿݃F���Y�^��/��<Ҍ#sW���2K	y�S�脘�+� �~z����AP��n�"������H���5��̗�����yif�Y���ǐ�ʠ4���7��,=�4[���6�m�j���|h��S��Է;9RH���/��.��;���	�z)� �c����zˍ�O,(�=YΨ�Q~���TQ�Zj���H�lqR.���IU���{R&�O���.ekƵ��e�\!���	=�I�sg��E£��>?�J2S�HL�H�z S�Y�� H��{t�OP]�Iu#�a�[�I3���r�����ϳ\ Ҫ�`O5C]�WG�hQQ��Ƙ��	��Q���Y�*�;��s^�� �+l�L�Y<c�&����O#� �N��1��=�5����e�]�M�ǠJ�D�8J8����vhx�XB4"4���+��M��]����б|�~�i��������Ch���5)d�ό�U@���sMi3Pn����\k�"�έ6	r�����UJ��н-�a��!��Ol�s7#9�~��\s��n��]v)�������O"T2�A-�6��n�:���.�'����kx���o��Q��::��i�wӘ>� qr,�� Lf�Z� ��"�gX%paW6��a��Ґs!�xy��4\���]�ݚ��=.��cYc�����#V=�c��3��u��2,2Q|Z�u�T�E��X��k��/�q�v$%5��3���7�.� �\�WH��b3|�323Ư�|� ��rRWK��s]І?�p�������pCPiwXԫ�����Z�I�Ӿ*�V/S����X��li^���
J���\Y�ۘ`����)����K�ܔ�kb�&��|�o�b.�x͘V�t���	�%2����>Go�����6�|�"W���k5�Yn�,?F��Lp��	Grc��n���K`�_P��qͶp�*�h��U"֧H{���p�N�:��	�M�t�S�&H���kGԒC���ۂ��ꋙ�J�7���kC�0�r�eծr[��Q<?��K|��VpЈhv�H��|�Cʋ����� ������G�������e�[�.��\"�R;ʉ-vI���A�;��dj�����H���{(B��Iz���������*���]�O��V�]��V��N���j�g�u(y�o��2,�I��^�<��Q�rN��!(wf��j�κ�_)�/��)����;����"�&.����U��'YY8�r��;���7@��=ml���!P�+����:�O����0.�
���dfD����:cf��/�)����|A1�4�<_n��p��Q�U�უ�&o�>[����j^nɳ���6
�p�p�4�p��/��j׽�ǘFF
�+�P�6����o�$�pJ?�w=��=)���M���ތ�ƴ�Iʋ��?�\mq�G�P�re<"M*3j��m��U�ԙ�o��)��̀��zE�]ˋ����=�3q��d��z3�j�-$����W�"p�RљR��`�v���dP�T�Q�(
+Х[�L�UΑ���$	uF�I	w|�]Zޙ��.o^����kη�@�'�z��5�4�٠$�t�yI6؈�4���pD�z&���	r�t|��4���[���F�W2�W�����\��"H
���!Gz1j X����卤!}�F�l�C�McA�<߃�)�R���/ou@���g�����)FB�s=PptOg�Qs	���E�!���)~y�§�%�-���*>IT4o�b�ˁ�g옿�{��EX���qr����=j��M�h[��o
����2Te@S*�G			��R���l����6B�l��
xm�G%�V�P*���fI�"6���p�8�/����"eo� �򈼹��w����nN�+��:8+ae�9�vf���+���k����7>p�̎�i�����y�����Vj�Z�S9�J�PK��j)�t�x�GO��oOp
�=�|L�4MM \Ɓ���Y�@��O��dO�O߄�4�ݾ
�R�0]ӕq,�ȹ��-cRK�W�=ֽ��͎|��]	�5ߩ���7nn��u���o�1�Z~j0'E[q�M����*f��am���4�4��!���.c�F]w��d3��uI�� �^�5V"�$Ï1m�_6 �L3��HLh�Ϡ��Q�ą�qԨC�cmT�0I���(���uT�'���Y�h� .�ec�#��1�}^��-Q���\�S��/8�\Pkb1��'��	c�Mdu��S��(��<�R��J�6?7.6m_��c`�xf!p�,Q��0K9%Y#���һ{c�sq�e��	�~�@���(�����NC%N�Fi\;kd�i�T�i�g����礤o��ȷB�Lr#�Y�;�4#�y�M�V���/�t��J"_�	ꕭ�������[pVLd�b$�+���wl��V�����K>)��,�"���4��$�����-u���2�(9���ʥ[�����w7��͂�n},8����r�僔`�_`��G��DP5UL �	7�G�D����;������U�z�Z�y��� �e��Dn�#%l�EW��p�烙V����c{O��}��݇{�����R8�3�F��8^��v�;����uI��_��z������I7M$���R�KHڒ;�������[����ʼ��l�¢��П��w$H��^���u7�k͉C�R�+�v��f)��q}EW�W�p��g��SO�Sy���ǵ�Ē G��@Ra2�v�J����(-+�bB����w~J�����mG���������{]�?�1;��W#�=L�����Ew����ws�@�]�i�WC�"�*rXF{�b,��,;U�E�Gj���Vn����6T��������	Ibo����ի?���j0>���"3g��[����,�.Em���	uX�����Ĭ���|xr	���EW�/'�4S�ԁkl`�7 �	
�w@�*ڪV�JT�!�����L������������ɾ��H�g���e+�D��:��U�d� p	g�!��Mh�H���Kpd��,4��-��f����&��<��坴��$�/&���4��y�ٓS,h���9F�r$~�]c�Z�nz_4�Ą�A�C`��J� �gOcn3�~=��r���I�\AʣFv�Z8/��#ó܋Z���nj7X�n͈z�����rvydxABf�wn���J4�Z�`v�H�I3mPLB �4��<�9rmxqmּ�*��Z�5�!���a@�˵��tʖ�|�-�,f��`��?��^F�0����I�Z�n��� ���φc3V��?�9�W��w�r^�cv�Ո�?�OF�2�m��#Z�|w�z%��xI�����e��o��Z`U��>~�c``\�5���W��ԏ'W������7�����~�j_�>�q��"�a�D�!��#���06��q9L�n�8�
�b�X٭��}{U�5�l�R}+
Č*�Lv��h{�\����mR��+�=�w�?�}#���z9�k?������8[�k�����
OUœ�+��n5��}OT��X�G��	m�y�s�GP�j��9(�
�����qoШ~�]�֣�1�p�������'Ez<M����]u��S6������[��l�͒�ӛ�������{�F�(�-d�c�WK��F(J�׶�V�^N�{Or��V���'���^�����w�8��jZ�o[�_���q[s 
���M�0e�4]�f���:H�h>�S��g�]M��規�4�8�J2��ȅ>L�o�_R����("]�*2B}%&oM��W���~W���;i ��!���,���-L!�[��R�{��XJH�6����.'�䓚qI�xG>�n����XU�:ؕ!N&�Gbu�B�FɟIM5:N��ҊGs�U5��lM�� RDf:�rҍ�����	�V7hc�
�8�E[�ix���I͚+^'dy�[�3w�
\Cp�b��)�Ш[�E�G��m�c{R���U�^< ���U�|(U��t����N�\�q.�
#E~z��-_A%PH_W�ߋ�Ab|q��N7�)�Y����8K�a���|]0��"��,��;�Z���$�9�x\H;����3��X��.&��zY���4-��ݚp�C%X~��Q_
��-���'34}���zY+�ԥ������4���g�By�D(; �1�LH!��Y���h��1��?!��_Y�'�e���d�D*$g������f'D��9>��|-��B�:�4��i�a(��A(Z�*ɽX�C�
�g��b��bs[�Da�D��4-1�lé����Fh㗶��i����A�2�ٵ�]�0��z6�1�皔K�\)#ܗLm�iD�,�=��ȡ�<�(��P�� R��4�S�y&�9��x��o��)�M�q�6�qiI��N��w=��}<W�tQ6L�I_�%��j\ko�݀e������Gڂ����gmC}v�U/d ��[��(�Pa8�排Y�����	��^}��?�mO�К$ ヺ'��E���v� ?��΂��b�p&�;�=^Iһ��H���5���Ӵѻ�z�Tp�y�U�ݐ��NQ���� }�!���\n�䞟x�IE��+(�$��Yv��
Ƭ�
�<V��V�Ľw�ު��iߕZ�Ny��P�4��L��vBYP��<Q�i�ҽ�d[��Q2��o����[�w,� �Xں�p�����t�x��0�WIz��U��������;�:��ř�; �ġz=ToPK*Dқ;	(r�)��7�Q�	߰}�e����w���(J�����O�F���i
�Aٽ��+��!pԊ�	��6�w���O`'�'�r�=�^p_٪��j�`Г����8�1k ��e�Vg A�y���wy����nbh�n<,3�@���༷�頗`'���]�p�[�9��pʌ�黏�0R��訍�8>gr�J�|��\�mޗM�r�����'%c�Nwӱ�����tJ�w�>^:�h��nF�0{�cХqa�� �5S���
��E�*�k	{�����L�x{�v���P�
�(
CEB��AT8@ΤW�"J�B����X��/��bf�%��i����]�35N�� ٞf�:
��\T.�!{�H���/�,�H��#�е���fm�T�R��/�`wcJK����5�rG�n��6<�����5��U���W�w���3L��$�uP"�%�^���^�Dܹ����J�E7|�ㄡkǚ� ���;���q�b��9��u�s�s,��'�Y�f[��Lq��pc���N���8j��`��4��B\5;#Zj�ɠ����7� a��J��A��(��������md�Ǘ�b�XYh�F	���N��Gh�,ZSje��i���؜Բ�C����+�4�}�%�r�<|x"��عE����8�>hc��?�OG� �/]1�>�3M��FV��N>Pn�sp��F��N�a�J���m�Ùc��R�g�l�R��0̍R���Y���܈�ݬ�`~�GIT.?L5��wF��!�f�"� }�
^ bg�/F\/`#��cغ��1(���N.7�АM������:v~�)Ow,F'�o
`W*�t2=]��*�8���(���x�V�tq����#������Bo]�]f�"o/	q��F�����an�D���n�yC�s�;D�6��L�W¿0M��3K�U��E �KDn��@d�bg�g��6+>��?U��y�})�{n��qa��ii�,��(���ω�q�g*;�x�|9$�䤺��R�����MG`IH�)��|�g}����<�6.ai�+3
9�^�y�X{ng�끄�s3j�E.;����)*Ѕ/%�u�]~���ݩB�I�g2@%`�N�?X��Ў�M��������p�D5T� ���>����(P�+�l��^ң@�^�*6�;Z*Y�J�\ +S��^Q����m�ng�U�l�iY"xi�U��Ie�Eo�"��bo��P�	󣘓�(���D,�;�|��w�lA)�%���ǎ4��:���o��mvl#�����ŉ��<�
�oG޳�G���`̹Rݵ��}�o�a�.S�y�K�}� �W�AZ6SӁ7_w#��H��E����&]�/��>7
��J�8������h����c�t��;`�~���-.��[�h��T!8��򧖑4�nm�П��e&$ �ԍ؇n�E�ѵУlx��Y �PV�h�슒7K<���t�p����N��,�{U�]���<7�>������?:Ɨ��u�Ԍ\���������|՞-����6D�xMG��q(Ђ$0ltw���s���c	�,h;��,Gul���u�>L=2ί������|�݄���{P�~�mׁQ�}6٦|>���6�s�7N�GC~�[�p
ʃ�����@�_ө-,z�����v���@ Q�p��Hn�{�u��<�v�PbQ	{-Qu�Y�C;]����q�}��`���1�B���;�m����^�Ѐ�5��ܼ�"
V7,c9���V���!ɩY��HD D�ߛ��ڣ��)�S"�
)_1������s
��`G�~��e|d�x��k�G0�|v(�4c��C�g�8�
�^�߼����DU�ַ�J���:�}7k��Ӱ˗�D���rI��V鐋�$8�՘������N��us!�޸�y���o$,#�E�h-�uS���Ŕ9����O�K�A\�S�ʖ��#<���������]�D�1�x�[`0�b����UK,��dҚ����(�J���P���o	�w�_HzD�^/�*,�J��o���u������r��W`
ʿ���L~�,	T~=9�2��f ����+-��I5��u��������X%����J��[�z��s����%	�%k:��GY�'���4�w7G��g�[��̳�&mU!�cDR:p����: kq�;�"a����<)S¢�ȭ*$-:&�L�7_�� �W�f�5;�g�l���?���t�/���h��NU�EY3�`���[f'q��B!�dl��*+� �������N�vmp���?٬&�s*�?уniOP�3?#�
L�E;���mfd�����"��T�2�j�s&������<K�hA����jz�(���:g���ӂ�-^>3) �ZӨ�u��4�l��<�X�����f���e�?��>M̵�_D��F5;{Ny�J�Lsʈ#�jI���>Y�,�Gܜ�������i`$�V	�h�U=��w�m�{ �7�ygY4Q�@�9#�u���N(x<��MB���;��̿L��+��X���F����;��:xhhh�D�RUx\�(��(��NF�i[�����(,�{�%/�&����Xm^����m�|�}i���N^��&�ü��f�"�܉���	A���վ8y>E��<.��PI�&�4X�Ŏ�s�B�������t��|�;�?��(�^���mK����_��\|������-����%�H��Q��w��3Z�������_V#0�@ :@U25-_f��&���}��$O:�@�� e�ޑ�2��{�\^���]q����$����0��E�Đ �f3_��gj���G8|f�a�0Ma�`�Z��f�L�D��o�&�1�
��B!����:ϑ71r�t�6�����ڬ<Y��eϩ�{�1Z,��z�S���n���ڒ^�1G����0-�!�� n�k��F\G$����·"�Q�nn�8�ȃ��}}_�� ��w���+�J�d������k��8\�#�%lz(����P�h�ky_M��C�ݤk��v �*����"�U�A  ��>j��o-��� !���6���f��##��":ႀ�@g�!��	$�}2k��)��`�|�°�s��ژ�o7���)Bn�~����ķ�+j��l1��M6${�ȋr��^]��.6c��|��M����?g�6�~/H/\����B¸t�W'N��C��d�`�	�G>r��>{�-���O��b��/Cxck��hE��ฺ8��؋d�`��gI�BRƤX�2ixHN��e�=�X�!m4���[��_'����y��A�{�׶����kޖd�P�Y֝���L���Ay�f5��W���VF��W�'�'��:�gvd�˓����L�N%��V�2t
�)6tI챏����
�ߚm��Bň%�Zil�i���$�?�K�[{g/`?�
/�#I,}�}3�N̋�jc�VZ]� 	
U4;ձ���f����*���LǤ��~���w2����$���8n�fC+L�p��`����ű����\sB�3>-��UϤ��'`�냵T��7�tu
��/>W��Xf�g�ѹiFR+8��_Y�E/�aD�FQ@_'�'|�I��H������F}��h��8<@G���$�A�8�]�-��N��j�lRl՞�}]�Z5�i��o8r]��V|P���t��%N��� ^,��p�Q��(H�\�B�ᮭ��f~z�Q������c�����@�n
�1xr[��E:�K��E}�i*b;��Tl;[���Ge��V[��[���m�Q|E��	Ę�4��L���k�D
���/�u���7��}RqcQy(`�.��/P�+:�����O�2��,צ%�f뀿z��+��24��S��v4W�2��'ʵ��}��<�:�-:F�Q���G�QX��iaKuE��"�����霜�؟�։��7I��`����D ������'�6�[cae�F�(�W�:J�&NpL!�P�{uJ�d^����DE�d�:ԫ)��S�@\c�l�4��O�7Z�(a˫<��u�cj4�?��7�P����Y�F7������zUS�X�q����R�
KD��u)�j-�g���+��@-	6Zos�S0�:Zxy'Ts9�ꑢ��rH�F������v��)[�g:�kl���'�~q�§h��;qi�F�~��J��E~K��D�E����-�%�:Fkr�ʶX'��V�<��/E�o�?�#�咾p�}
e�G#

^�,��ϴ��W~�{-_������sɶ^ �K��H]0���V�
����1�6�Gן�h��/ά�xFKP�^�H:{�oXlxVHYEB    964e    1150R�]�	�D%������_b�Tؑ=���3U�^��{Uc�|3W���_���(?z�@��B�����j*o�� �k�<�y�cG^F��`)��k2u?��k�&+���5�=JřZ+�_���ҝ��FX����s�B,�$G�Ĕzn�,���`�4�K$�C�Ev�|ڋ�n6�KE��y��mw�������36�H�^xasZbj�7ң+ă�]HV'K'e�
&�>�B��P�e%��V��r)��
��pإJ\�Lԑ��	�I�δX��뺛1��+����κ�����+,�MuY�nˉ��-��J5dfJQ���<�&����{�)�o���C���![�_����ɱY�����q�-���B.��ʷV��J9��Rn��ÜU6�O �3M-DZz`�}(������FA� N0���r-�*�����-�Lҹ�L�q������XН�ߴ�FlT+�HCXOx�y)�Z˞0-���DP���f?�>}�񦿒Q�A���!-���Ɐ�M�S�<p����ωl�-���/!�����\��?|`i�/7�0o����((���$�41����U���?-�Xlg�*nasK�b�lP^�����v>��M���w:���~��[�����j�";�e��������]�4�wm�h�xg�����~�O������=зUMf���$z�T���/:ɞ$��=g�!_#Q:�{^A���=�^*qܾ��V��5O�e�w�s*�2��TLXB�\���
N^.R�^E�Qo{b���X���S|�������>d�2w{�cp0�%ｄ;�W ��u���%3���"K���/A�E���W�9]lp��+s�Z}M"�qh���W�SU�����S�E��wXiRm�����}�a��jDA���g��p����R@;�sBl���hdm��l�F����̂�Ah�(�ު��LE�V)�, ��&S7���L,�Dj�"Km��{��ho�Z�f4�l����3���ä���5#��BX�ȍ��F��~��^�u�2�Љ��Y�oo
Q3��	�(�l�1�EMc �D�������]\h}��ݔYd�c�z�?=h�vV��oe��=��I�י�~y ��s�G�C��Ύq&�v��Bģ^1zKNc��P �nb���4h�>���8�՘�a_�
(�E�e�Y���4ʶ��$��A3�#ŸL�}�?t�}��8��^|��Qș��/J���ߚ��y9r`����4kX�fЦP�sF&�z)�H�ez�l����g�;�	����G��n�����o�e
$<V'HFE�H���L��|�Udu|�&��j�_4]�� �mPkRR��8�8�{��ĉI�v�A!�l}��I�~�F�C��s{�J'���Ă��%����,�	cdr�m;O����AO��Lc��h�M��2u%L߅('5p���: ���q���z1t�MJ���"|;sBL��>n�(�4��@�k�i���-�J7G�R�����O f�ESGJ������o�9/rBRN��.�Ӂ�V�}p5��3	;8����,�(�}�=��C�7�����#����(R�8=�k�A@���j�֥�CB�5?��{��=[����.lٶ7���J��}��b���.4���*P/K��lx�zLUN�8ӳ\7����u	�nŴ���d�����Gw+=����$H�Y�V�u}��U��^��NcB��wnB��}d��E�8��*�b���)���5�e>+#6E~��FJZo���(/"�@ݯ������ 71�~Ca�UMw�Ï���~"Bg��&����t�WJ!�'X6RS볣�Ԛ
����p+��w�E�W@3~.��Tl�D��� ��R�E�f�壟U�X�0�̋��n��t[�~�`~*�
d!��Z��J}��/51I����4�^���@g~�}qf��_�_l�lT$�:�|�\�(��7|�/_ ߕ����_�f�?O����l�х6�j$5��n�_��tK�iz�����f��|�,�p�I6����,����u���Ŧ���ו|wA 9�G�7V�P|�}��F	����a=㙀��ᜆWg�ύ���3�{���į�n�b�}��ݼw��f���]c$&t������~��2�s���=�eԗl���;#��n�Wm�*�"{Wc%���$��m����p�2����s���Wwq�*�öO0�q��a����d����[+�$c�����{f0������Ѩ}�{�4	�)d�����97aO^Gr�µ���a#��
�a��A����U�X�<�6@P����F��T�	��>���Qḧk&�{浍���5{~N(�ό]ځ�v���B���Z�R�����[��!YBf��k=�za �O.�	��|KG�L�4��J������f88�Vk�u�w��Z.��f�:�.��n,˨!#�Z����Y)�/37��NЬ��j��4{��<@W��Av���g��m���`W��qy�)%I= {���M���	ߢ,��3�Qj@J�0�b�	�`.�+�6o�G	�ɤƼ��lHb�
��+�K�0P��m��s��g	/'�FZ#c�<$U�|�{?�����o!�����Ѥ,��@�e�鲸���R���t�ٯ��>s0V�K�q#	�{�5��Q�fb��ulL���cO��e�J�G.ˆT�2'� Ȑ3���֡?��B���Շ !	jX�je�P	�7�vD�*W��f�R�wa��G������"���d�P��Lj'����:�FU���5fc�$�L�>n��d+ ��|���2�"c.2�^��M���GFj�"����l�t!�y� B�;�o�(G�#b��>7/�߉<�g�ˏ��:�GP�b}�JZv�Σ��.j[~}l�:W�J}����A�f�XeEHO�J�a��3���$�ݽ�x�Z@����M1����" �&����)��#�GA*�գ���!t5.Δ�G�=�<���S�B��^��+� m���q���&���6�i��8t�%��q��~J�<�j*�!����Xa־��%F�����d��bƍ��ͅ�̶��X������cu4P�}���ߖ�^�l��f�l��I�vy[0߂�Epw��zI��/���{���5�*�@OU����Г�A��9�����ϒ��߯>�w:�wFH��ZWq)���.1/���),Y� �q����1ۥC7�!�W���	4��͒�zAG���:���E��i������`�\�W̑�kL�(�C�!���7$>^�r�"v�)u�mࠖ:_��$TYq��H��sWݤ�����Y��������&B��S�5\"��"�f|���Lk1,K��8�`�n����MӃ��V�$'^���wަ�KU1X�y�uV�����9oJ�-����M�\��1�s����r67��H���4 п�fx��謸?x�,�%5�6Ew! }z=AJ�9�"�=m�$��O9�P�=��<��\� ���`��Tp�l���lO����hse�CR� Vn�Q��TUo�댽0ׁKD+Q ��@G������=�Z�܋i�FR��*��T�`�p���]�^JW�h<m�����#���� ����k��r�u�E���b��>�C��R�qT�����`�kr�4���N���"�p���џ�?�0���Tƫj|�v_�����>w�_�����`wX_��������n9�A��B]���~4 �3��L��t�O�5��:�[�s'"�����:��}�{a�}�9��m��AD�6,�6��Ҷ�4 nȺ�_s�J�w����9�-�|����Q3��^pd���A����)�­��m!@�@����T�$i<�n��6!7Y�g��G��,���@��/Q���n[oN�����>�#%��М6����u�@k8׿�Y�ZZd2�ֶ��[��k�c�&ǨyC$�YX��m�D	`&���ZSqiq3����gO8��6򾒗\�D�ػ������N%�5ɲ�}WO�Q�QӅ�t��ďs��H@:lR��v ����=A��`����Џ�F4g�Z$���(x��W�%`�{��w��7�/ r�8����&2xIoo��&����]uЂ,D�j��3�+0�N��dK_=>-eI�����%.O�>�(�Т�����+�`{+���Q��;�nM9�Y��ݶ�n�qSo�]q��(.�\6��9�D)*/�{���z���W'h4IU�5/��X�^�#�ۤ�i6ƽ� ��fM�ZK1(��Xn.zI�^�#L9���=�V*����0z�&Ec��0���aŻp!�Vw+��\TO-