XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1�q�~:�n���I� :�tt�?!E�.t��W�.�]#ղ�U��;�ߴ�*��9��c�R=]��Z��.���W�O5�h�܄����(�°+�g�I��9<��	���l_�}Ҍ��NY��� ln�"�"vWC��b�ά(N�gw���F�'�o�D���g9-Tz�?�`7��'��������Q��L��ц1E�6(��NZ	?�\(֢ 4̑�pd�}�V���f�s�h���%&�o3����mR�ޱ��C�긑%p8�Յ��鷿'�@e�E���-hG��?�*Q�S��h���I��}�������F�u�3l�0���'WE��?f�ΰ�˅��-���J��N*���	�D��zB�nȟ�eo�T"߹�Z�*���������V���q������p؝y�A `�M)���*�P�x�̓����s�>�qk��ߚ�J_N)9����A�!p<����� 7w/�mQts`��]�A/�僢�7��4��e��s�4N���T�q�2��\����:m/;s�aC�_��/����	�Sq�<�5i��c7��-#������b�zn�.�ɇ�7ڰ�e�t�6�
z17�Ý�Ȱ�ՙ��p{=B�t~�sp�&��Ń��Dzr��ʥ�b+8{��K;��0���R��NGg���o�+^���f}+�|�H���3B�!�����׊v��c8~y��
��6�z"����q%?w��c�̻1Lnǀ�U3:HT��K/XlxVHYEB    1427     840�ux��a��� �G����r�n#����=�v���uTG���o��k`R"�ǎ7S+ڧ�~<�CS������T�ѯ�$�Wv��2x� �+7]�n�y���e,At�(I>��MФ�����Y]���f�?�\��{���8�)�]"&�=�0�	xj�u7��Exډ,��8��B��詫e�4b/�Z���Tx� ��d���*�L��*C�[��p��ݢ��F��ڳ��!}+� G��>":�E?���*�u)���ā�{�Š+׹|n��;$�u�����9���8y��?���޻s�uۡ�U�1'�&ʏc��,�l�]�؋e*�>�,���S	�z�L�p�7H�� W=Q���6xlK�s�ՠ�S+TN�v_�4��2i�*�.d�В������`ԓQ��1!�#��P�b�4����cC��'�+��g���8�-;Z�g*#(�
��gj��8Z��9���;�C͉#�E�2��!���5�$����Ύ��US� ��!	�`v��S7������c�;�9⨍r�O���1^K�E���(7}׈o�L]s䝗�%t(c	d�Ӡ���P]zL��	�5�*i��	RZ.��H�6 �ᥩX&�y����/�M�s��߸���9�!�?�����9���IL�R*2�T�b!�-�L�Z˱���6#oKI��)g������lJ��}?����5�juӄL���"����k���gIÂ��b���x���|[�-�A�N彔r[;Xk�P�����u5L�0�	�YF���P��8�Ng-9�42e��^�X9?XH�!0i	������q��*S�������k����=c]l"�ᆿK\�����BB�0���ǥM��jlƹ*A��k�hh�4ѻ��J��I��D� 8��}�^��N��\�i�.:�{�����i>�2*���R4�L4��*��>!(���0���W�9����U�f	��_�r�Kk��6��ɢT��'\��O���uY�o}#� 	�:Y ���v��fco��Ȗ+��$��ˊ!�G�S���ʰ��n��2�դʰ�>�]N��c�`����ذ%�Хy �:��gn�f~�r�I6|+MB�b��le�z�)������q\R����u�s$�^���
~-H\x~E� �zz�;�.]LwJ>>Z�������D����#��S8�����e�"���v?6�:ܻ:TI鸏�#��̢1m�����H��_C�Pf��{�yhd�4�y���ˏ���� d<��Jܰ�4��Y��u:~��]n�\��:��7Ny7�{1Na"�z�׶@�̴�0�t��ܻቑ����q�S�Y���{U&���8�@?�S�Z�s�߽�YWpSɜ|���zu#9�Љ`ݤ�9���q�h�Y+�F��� fw��a�AN��߆ٜ//���pB��.�k}��k��W`d�������]�|&����X|�	ݡ%=rEi�2&��6�6��3������a�|���ceܝ���Sg�P�հ���t�y��S�|M��,T�Z[gxoq�F^^)��R�!���0g��w��C�B��$�S���:e�_6c'
2��l�P(~}�׷�}�\
L��k���H<g���������Gͭ��ӳ��h,�M@@P~
Vёu4 �s'w?9��+��SƝU]4��X<�1o�$��91i��:%�9��� ��C/'Oѽ���k<�R�0�Yˠ�P�{�'Zd�B���TaY� e�)�0�w��	0� ��scj�p��U���?��<�n�����5�Z̛ξN���\�qO(�>z�(z�u�rm�O�r�ǒ�ώ��H�Ҝ+��\�u���FCcB8�F��B�0�;g��{�*�>t�9fxD����Yr����g����4�Єֹ��b�ov�6�����R�W�n�m��~�+`E�Yūk�7��W7r��2E��_5M��p
�[��|%ߐ{��U�J;g7sͺ�b�z�M���xX��j�&I�xnL�ݛe��V�(�;ِ�U��u!iV-Ea��