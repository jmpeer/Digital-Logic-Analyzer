XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y�{v��?'N�������%Wu�Mbv�����[`Y�G�oE�����m1$�+Y��)����W� ~��E�-��Fr����@Ld�� ���9��O�κ b`�%��3 ��}z�k�����g���b�e��]��YK�a=eG��0��?��vj�D@[�7ġ�6;ya?��&F|mbs��/o��]k_�2���=�@Mbm�ψ>^���p5Jy���h��CJ���޵������=ܫ�_!}�E^M��A�B�r�$�h̷��Z����;E!���]\R���Y�s^�	T��o�O#ӡ�������`�"eu�c�	�N֓a{��q��6]?�פr�`�z��K��B��M�
Q�{��{OCB e�d]Nv�lu�z���(i����=V�e�|����O2����!0+�V�N��y�ܿ" '�Kܯ���9# !%�}wC�[����2��h�<0+���d֧�P>A���կ/ޞ�/x$̷�NϹ߃6���f�<��;�l�cu$B�!�G�WYi@6�*����]��-�w�Ngԙ�K�/e�@(������{4����m��Z�~���]'�xO�q�������]V�,����Y2���:�;}�\'�/l|�W�l�e��z���2c�}]��"%j3C�Y+��Z�a��5��԰P�*�&�D���n�I�Y��{��&������m����cƣ���|��͂��;����mXlxVHYEB    162c     850�K;��{y��}W��X�f��&ڙPT�A�ו��R �-ZV��j�C��v\�va�|y�z���r#=r4TLyIX9P955а����e�d����x(�E��3�CB�λ�J}Z���¹_�Z|�U�Y�:PI��|R�0#�zb�/�*|�9��xb��p�r�O���?�`4盧\pɠpey�U`�+���r�X`k5�W��{eX��8lͼ^e�7�Ț��]�(,���4����	�x����R���Kq���j��U��M��.p��"w���u�7�֖3,��7��"�`>�emm�	���P�<>��(�EL��g\�;��&Ƿ����6�*�E�'���Ƞh]��*�[-���30�lq�B<�T�Cf�	��;*p	]��(��%B��-���=����`����7L���K�/=>�r��ӮX�#�PU_=Q���EC<������:��s"p?Z签K j��BҴ��_�Y��n|��s����t��>�(P*'�+kJw���!�����ٍ��㮊�����C�'��H|�;0�3�{5��kP8�A�Jc��.�#�h�MO�C��Hk���4G薺�����=���y��G\���3W`ʓ��A���d���CxEI'k�v�Ѭ�6�,Ѣ��פ��q�<���������dsGX�?p��.:n ���ah��ȥ:'� �dLh`ҩ�47��C$U�7�ZbX�UJ��Z!`�����+�C^�x[A@�$i)Zo��+_���ʙb����_�d�"��
Zw$S��A�U9�✽�����������)�>f%�댒7�﯍	hUK1��G��\��k)�-����L�>*$�R_ߠ���x�(s/�9V��1ql��ܧ��9跅q˙fE��f�/[vàP�f�v�w�<��Cp��� ��B���8/*�+	��E�������!i�)�US*]=�x?<g�O��I�¥)s�e��7����ydeU9��H~B��h�յ�ы�3Ѻ��
H�@�p�v�D4�����}a ���Ah$��$7��I�z��b�A��5׺�Y)�WN����v5*�¾��:��X����/����	̡̲;�=����BO��$Yjq�?�7�*�3Ј�-9�Ҡ�F�[�d�@��`x���h5$����![l����<Z���8��^%QK֕G���TV��aa�zm�Ut5)�C�]�4�t��OW��m}w�_�9�ඞ�f&��I�Jb��k�K�hs��S	·��HqjS�.p�b�ռ/�{4d�'�7��-޺�x,B����)�ff2�AsU[fe�n7F�T)uc��ئ��f���W3��9|�~[��_���u�2�����)��W��R{����U,� �%"M�]�������t0�;�Fľ�)���f����N�ݐ���˷��;�|ͮ���VCU(Y	@�� �}�	 G��봶Eed�}���sO�׎[$1���C��w��*��!u'���0ۖ����k5�1��h�.�i�K��P��ǳ����@fgt��g_��N�A��\w��m`����hY�&���]Mf�=tA%������U�w��Z��DY�HLt���̔���y�����X/V�x;�ޱՌ�flg��2e��q���D�2fq܅]-�)�����?Tk�g��4�i���$ ��TѮ\x�YZ9���U�/t�����d�}k\�5�gP15.�%�� Y��kB9u~��n�I�.����P��cj7:O�I0��x���rE�M;w�,��vￖ�s���6�Sʜ�{%�d�,�H���E�ǫ��cc͢h2�o�v.�k�Q�>Y#���q�i��ʐ�����'a;/]���#%��	�
��6_��/�P��uPvA� %�m�W�+�r���QQf��-aȳJT�ᛟ��M��u�j)@b8��'��P]n䓩�uh�2[�/ L����7�����?l�.磺����R�
@)�/_���OK�RZi��v���;�JI�_��K�f%����Vy��	p��<�������'����2�G���M�.��