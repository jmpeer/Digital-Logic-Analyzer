XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����&Ue�<�U�=���B�I	��_H��(��^<�9�P�J�xx�����kLb��[ǣ*?��T���@��Sf��_�V-�y��J��L��8|J�j��߭�L��-�[���۹�|��ND��ji����M���i�Z
UP�m���=՝�.L���Մ����ԤW;X�k-�=]�$�y_x(*�R˥��AQ�T�ΘDD�5��L�@ �xo�bO�D�R0,+)�g]�_yG�w]	4:}P��\�����ӣ�.��t��G���샙0��:�톐KF�4]�!lX�n$$��R�>��錸aV�o�v�fϭ�F� N�M�Hb;��{��ۨ���5g�X���@�"�*�u�a�������c�hl�j��{x�MR��H�m����L�C�~�9"r %�KsԎ�ֱ��`sZ��E�"�z�u�gp�ۚPL+x���w��鹤P0���<CL���F��7�\?�<ϨcD��N�����n]Zi�.����
T��r����1݇��.�K󯎯Ã?류���IT��K��Av�fܽFf��Y��F��.k%�+Y�
CAJR	f�c�.�\Odnsp��ʦ+֣6�|O�AL�O��-�L��l�V]P)�x��˯�u����6���_���Ju���C��2np�Ǿ���W�ň&x|�V	�R"��J�_1K��14�����h|���wj
Ŏ.��'}j?�o���UW�-�Y5;\y�)�v���K��]{XlxVHYEB    7744    1780"��'���5S@}|(���?u"���:V ����yמ���g�Y�4R�O��� �)��'��a�0�س m��AX��=�eK�/�d]A��ڗ���������M����I����I�䍮MK(*EvA�L)��t�_�S犫C����	���;��~-��D�	�N�O�$�Jw�$��ʩ�`���XK��K�������j����	��f��_����+h�Х?f"�<����O7�o�>�1���P�����=�\�IX�|���糢�>Y�>W���Un�:�m*.�R4��w���աG��]���C.V������}<�L���5�Q|dS��58�i5���7�^6�߼A�[���a�Y$�1���D�rp�(�ׅ�n�����d3��D�i0�5��c����c��.��6�$��՚nT��~�+_����\j}43��ڻ��E��*;�1Y�圛#���`���L�!G5��A'�7��U���sj??m¶� 	�2��k,�d�/!��{O�'N�n��C�� ��� a���'�{�CY��km��t����]t�ʈϥ���0��/
pq���d$P�nt�@Ԣ[��Y�NQ"�t�~�*Wp��{M��%ٮ�֙NT�Q<y��G���:O
�`v�Z;�(�i���C�s�?�9~��`�|�𱝽��p��Syv�i�����ۡP]7.�� ��0��N,|f�=�S3�G��
��̌:CV2ek�	����e�ٓ��!;t�Q�h�#���:;,�lI]��X�tOH��21����N�w��|��l�D�i-(K�_ǴX��=�34��G��`�贴.�8q��5S7_��1nP��8�g9V#�����[��hi���-!�p�'�ȟ�ˁ����D�O�BP�_0n�a>|��B[�7F�<i�95=�5q���m�t{K|i�ViMԞd�P�Kд��v�\��2���D�L�� ��B#=[[���U�AQ�9���v�Z<��	�sG�]�3�K_u�[n��f�ۍ5�"�M;5���:E�~{�N2V9�S>��\ny$v�< j��<�n�Z;�}�d*�����.
/�ʵ]�o�������a�K^&,��d���z�y���4,kڲ��FP����@��RPWC�\3-��6�.(�r-ҧ���ha�F�����w8$NF�:��NL;Nr���$�9�`�4�̮Jr[��"��:<��:9��_�n� D�m�\v�&�!�Ըuw�U�����&���Ҧ�smN��t�j�D�/W��0���N�`sr�b��bL"Kz����z^gi&��rJXk��d�:�|:5J ���p}�i"�$����Gˉ߻�6��z�{K �/�Vw����م�T7��D���O0��o�m��-��5��Da͠���4 �~�K���I�$I��&�T���H�*��q�~��	�z�F|���R}'lI|o���N#���9�eذWu���9:^w�"�4��L`���K��	x�BEz>��7�~���z=��pW�n7��6W�T�Y��&���@=��I��vR��
���UÏe��r擥(�v���?u����t�[�''i?4�������M��b��=�\�ka��yD�Xd���	xη������E��Q���p��V�0.�k(� J5X�Cv$`鼏E�ğl�ˏ�Y	L}�G9XL�s&w�>�s�?�O�>K�����@�C��$�� z�G�<s��v�����50�����f}��� R�yG�P� R.n��.��|�)��@�p�gT��- #�v�3Լ%Z�������r�0�:@��U����>��r��@���B�����w��0wU�=`�:����	���?�n���yf�v/�k&⩋N�jcGc�4~J|Z�k�ӥq�m�ߪZ��S�4�.���5HWA���΢G6��|���<��-�p��~[��aPMB�ޙ'<�7J���2��_�{j5�!k��3'�8�rl����US>���E`���j��$�'�hLh��U&� Tk��C���!9�ώ6�6w.������P[rH�XG��B���l�2����0��K��Qd 8�f��U�2��Hx!��ʬ� @����>��_�}�ȸ��ʀ`T�ͱk<L(wmn,ڈ���AcZ|Gw���D*e������a�!	|Pm����G��騮#�D�4�N�����k�g���rd҇�.�z֯$�3�7��X+\�J�\�G��ch��Bƶ�|�wp�&���_R��PΪ�Ck�=Yj��3
�Q���Ŵ��bb�;�|�?|ӂh���	���I�RM�.��<���t%����/���>���?n�=@Q����5�c���^ ۇ�$��9u t���7T~�o��:xb�����]�M���I(��)��%������G*R����]T��>�M��a�v���|�I�^g#��[`.�	����fXN��k���ݒ��J��U��c�_X��'3sc�ĩ��hK��%8�-EZL�I�P̥�A��4���Rz߂�{$vI����&>E��uZ#��:�9��w��[W�� ��y�u�%(���@���*�ӄ�?lj�ï�Ȑ6=f�KIrfj�ߛ���p��c� �i⼳6�b@���Ý'�ֲ�|�ZYd����Qv!��o�K�#$�G㫯�\�x��&����uܶ1�l�axDj��4p�z^�YJq�r��d�˼�N��:���ۢ?	�FY��F�۷��^��H�Ybks1��'|߳��#R1�IN���r,{���lz���l,��5��/.�?G$S�<�Ą�2���KP��hD���a�Iq�>�y1�GR��Y;�g�K2g�߯FC;�]�;�	y�I��$��v����A�����q+���pՒ ��}$08�Y�|�c�����&�%QT|B����8ܗ���z��;�^��wxr�yI�d��)]�N��h5��[R�"�d����o@O�wN�u]V�!ÑE�{�>�������#Uc����L1n�+�����֒����'��8��]:\@�&w�k�fa��^���8�n/�?�M u�8"xG3��� ��hKѼ�l��&ֵ�ż�H����hĻ`ho��!O��完A��PO{���P�՘��z
"O:��J����;����@�z�91�]�Մ#N��֥'�	dG�HK��������@3�
X�2���ʈ�jcr�$M� ����8�iw�Ĩ�����E�͋(,��*��G�*�^��~�5v��4��mP��ta���{a��!G���Woô��)=�KM���L��7����`���%�a�JhW�^0ʰ�Dg�ή����T�bi SL7��9�%{�6�:��V|�Q�(/���E�_��H[!��
gm㝋��%�_��k���6ŋ��X��cÚA���4	��Pp������Ӑ^;ZP����w�r"��Z|�<2��F(r�0� &d���y݄*�جO8gzZ�9*C��?LI���ϧc�&�1�O����#�&c��#�/��P(��Y�R����ݲIԷ�k,x�z6L����5�{�ƩF��S�BͫiD��C��E��2$���o�+����),�����E�mk)j%�{^�c�o��?+RiѸ�����="<�o2���BNI|�=��7<F	��Ȑ��an��������$�4�U0��uM&��َ)|�����h��)	i�t���ˉ�������@5�C�Al͹L�%4;7fzgY�r��})lϮ�͸.�!��$�<}������H^u�$ă�k`��^��o�g=c��"@��h&���i��uȪ6. ��o�OQ�G�T��m(�'����h~�G�n/^)�<�4��zk|�UD&�i�u��p��z�с�nyh6\�^���Ѳ 0.☂�dXl��v����*B�V�O����W�~����GX�yp��yH�M��:���&�� �%�"�PB��Q�W����"l�(�[��\M�S�x�N�-�A��<������uZKi�{
��:s�s��a��A=~�a�1�=�|z+���
�*:E�(m�Δ$�8nK�3�L�(s� <����(��Om��&7%�O$@!0$F�,*d����X���/)Ȗ��*�|��|�E.��_\k�L��6����]g�6��z����%�R��9�� *�(40�c{qè¤��U�m߾����;�3&��!ŵ��c�q�����mv��c���/�S�{�U�M�8��X�1'���
�ۣX��?Jv�P�y�����W,���۾����\��K\G$'��y8����9�K?�B�2�\�|���B��E�1�0W�!3⸚����v!�;�T�х^d�mR)ў cî�!?�y��0۲Օ���1wdi_^�%NQ�܌�<�����.���ͮ���ORT��f�)��fi~m�v�z��h���s����W�l;|#�<gۏ�n�Ƙ�u�l`����S������
:b	��/��8����"'j��i���5^��[3�m|0����n�Q5H��%���]KM�z�B�[���&`�y��@�G�j%%ˇ�V�]`���T)������2�I~���M�CK���ΓL�ԅ4h� ��?��������&n�&8T��:�([��hs
mt@V�ޭw�~�-/��~��^�3����q��EHϥB�ހ1z�`��<VݼU�-�N	�e�Z̚=z���ag������FAU8HÜ �*g��UOH%��4}�)�zX������'�$E��G�����;/�{M	2������A1��Nm���okZ��{N�d��b�X�*���73ؘr�����K�������8��0M{�J���B)��#��˃0%�b#.�K���d����oЙ�P�i7���f��u�Iaa���?=U�F�선�k��c�5�u��FTa�<p�xP~N��3�4�$s�(�B[ܣ�ԇٔ�i)%���>� � k�,T�b�d(@�"``N�~�T!`�k�%��^x����+ĉf��@ڬ*��;�q��B�l���U'I$��(ko�A� T��F�_B��}��Ǝ�Uo�I���q3"|z4:�7آXR&>�	߹���9��i��f�l;	k��B2c�4���S5�ą�&���($�$��Ϛ�To�_թצ��>_�XW�X��ͫh�	G��������@vD��)��u):&ܓ���c�R��2$W� ���/���$>D��j�WB�L[$.�\z]����8����n-̣�~�)g�f��c�z�?c-���J-\77�J��JNO���dU13�nnO����1�	C)�%��2QFJ0���6��hl�AKb�q�)L�ɟ�����Sn��d�+�)��}�P.�y��RwA���Ӗe]ɹ[��5!ZUz-�-�;1|p��%��F�o<�T��S)\GP�s�<�%�p�/�.7�:��&whb�`�6h,�p/;*�����SRbV^���?�����`_����fu[QE�uO�� ������������6@���8~�Q����<�*�a�5��<ۥ��w�qP,�2�l���<�X��d.{W�_�9�}e��g�g0q{�Ѫ'D]\�^ W������r����1#�x��B�MGU�$gFK
!���[^.N�zP��-����Pʵ�����9��ªڲ�[[s���Տό��`�Gn�Y�����L�J�_�j4����F@�U����np*6��aqK��ZBc�cb��mc!5���1��2 ^��ξ?�E_N�Q֑?�N;):)*R��/>�8���=e�\WD�/���!��2�Jh|����D)��W)M�}��@��%<��Ș`�@,�*C�KƜ�>>�STh1�.tŒ���*8x���5Q�!�FܬTK]Ou