XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o��L�3���)��(2t�t����a8&\���?�v��9u�H��o�M���a�x�5���� ��bH�������C�I��~	 kqy�`_�Z
#n�xq��H[~v-@�ߖ)9�Ʋ�7BM�s��8^!�침k|&(0d�*T$��wh�O���s;����*ޚ����x$jvC�˹3B>]Ȕ)���J]�X�S_���~ء�~7U�������O���U$�ES�@���U��G��l��S�b�ux�k��L�AR�>]X|WwˌP��!�)
�O�G�yMw�zn@��B��:���זI`��)5�L�n��3��5��'5Wzc?,R�Y\��1q���YR�q��G-�V�O���%����Ꙁ�斯q�+'�r����4�|0o�7��iД���,�6U�WN�l�/ �l.�jZ�3��L1r�Xzٓ�)xG�]{3L�Ϊ�L)''�M��O���C@*�{�=�)l/-��z��*�idK`��O\��>��3Lc�D�)X�ŵ��dT���Z�$L�$�����2��î�}�0#j{AZ�Z�U����m�m���%����L��`�ƨw'���1a#�5��	�Dt�C�-}�	�De�����`��b�5��GOR�3�+��^�A��7�,.���6�ڹD��./O�JK�3^�����Jθ�WJM�ɥ�m��^;���M�T�0�`DW��D��aO�.��i� �9)�,|�Ȭ"�]�/Ư�S���O��!�m(�=�ilXlxVHYEB    29da     af0}��w�PJ뀋@R�Q��v~ҕ���^���\����_�ijW�H*[�0�[ ���;����S��p5S���z�^}�)���U�:Mu��pN���Ič���#oT���X����y	��o�#Z��Xb�! ���7�nB��B��\�];� �<wK;��E#,�n�4�t�-ɣ� ���P���n(�/�	�Ѡ�b�&��?�֟w��5���I��p�~��l��<�r���Gi�ŎԘ���]E#��W	O��6Rق,�$��㫩#UD����v��^���ruA�e��A@�A"�yC|��� ��W�xRE�Y! �؍:�Ϛn;O�Enla����a.�m���^��=��_@�Og[�a�6Z���Y��$N�լ�h��=�O}�
OOGOY�dN/f4��8��������R���'ׄWAO��EǨZ����5aN���
^tɤ��1�Z��\���n��x��S�E3���Γxw��7u�?k�т���ܺ�ױ��v��.��nФ�m��j�P��H���Rש����\l�e��DYrh,��輈���������{������Y,��U��d۩(Ań]��)��q�#� ^ȗ������s�M�C��yk�AF`�] d�Z
�k�5�C􉂽?
#�}�.V�h��}u݂�K�������T�u��i��!lvBh���1�3��}7G��<��V=��:O�ԝ��"��
�1Q'�����S�IYe͂�!`�'��X'u<�����G4(���W�@�����$���ny8a��I�Ξ� ���c�����7N>�t�X�;���pSk�2�E�����=��>ܱģH��;���D�iBN$�
h��wgM̍N���
B=�t�K0>~Z�h(�j���:o����r�:�6w��ڥ���3,�`�1@|�SҨ���-�M{;��f��ӵ�2
!��-�P�U��H�g��Ԗ�6d;���m�S��� E�ǁƪ�Y��~�?�s[�����e�gX�̣���G�j��w�b��r�������/��cr��(iTp&8C%�]�]�&uZ��j0��#ήŚ�yo}ٟ� `l$ �Tƚ�U'������O�;�u�H���! _7�ԝ��u��0u�
q.ʲ#S����p��ke�n܊;�[�jk���)M�@��;��wo��/���q�Uлkp��[^�(�s^h��8ڛ��3Fz�c=y�
�c�0dԪߍr]�艍����!������t�u�9|c�H����Jϡ"#���Ԧ992c1ˢ��*8k�\F�sS��8a��x$A�e%3B��N�B. {�Y"ۜ�%T}⊑��|u&�-���&���В�
��;dc�w�'&ykLټ0ϫ�������ѭ!��������@e'N	U��,c�Gp�.�H�9Gek\�}���-#s�1�1=�|��U���9��W��q���-h�Sh;�{!��>�](�fk��竤��H	vR�	�#�)���w�Ņ�/v/�x���\8b&}Q�_C���Q�!FE�Y��l�>$�f��y.B}62Z�򇺅Lt�O'�e���?6"#Kڽ9���K~�,��ޏ!�o�?����Yh�%Q�g���� �V�ev�+�n�u�УZ=^�M��Q�D�3��!�+�.l�*��HusV�-6���/���jqv��f��X�	c������6~��N-=��3؎ڙ0�Oh������I��5!��_3&?�W�%Nʏ�1�7�J-�������&}ՆHu�|Ϫ�V�S��	 g�������	8H0����aEzS�C�\[�a⑁_�����z��Z(��}iZI�>�e���!�=|XW�jѭ�D+ѕ����a("�젏}�����*��aV�6�}�)W�|���c���L1홸g:'�O˝���<�hW\���4�x"���e�۾�����U>�`��
r�����lѪ��|#T�!@�P��t#R��#7��t(X�)	A�xF��<���H����M���yGp/t4*�+��]�/B����Ve�	�QdM� ��_���ӄ��<n�aγ-xf ����S�9�j<��pJ�p����q��5n���W:��nVw���� ���k�Px>�����-ZU�Y��S �'��dFT��-�G��b�3PZ����z�R?;й�Ս���,��_ì�T�x��,�Dl��bE%��[�S��|5�*�8[�j�8��(�.0���0�r��Į&�,�9�06���)a�=Ge�ꍧ}��`G�0sO����8|/�B��!��-�oڡi��.��ig�?F��L�!�E��$k''�j�6�i����:5(�/E���ڶ������ĆJb���o_��`Y��15���y��D�kGJl�,R��L��er����zOp�y���JȾ��8�y���.}�+�X/�m��v
�`�_�R��J�}�V��E�k��OZ���Y��Ur:K���'���I'��% =�mve�~&�hD�G3�/��++���W��R��@���k���r��8��y�<�.�O�gO�,Ԏ���^�6���h�30���]��Z��2��:5
�L�Pr��W��ڷ��OS	%}3���On\*L�ï���b�VK�I��b���.'y(�hw����ԟb1��	�4t��#�g����J7�_V�G�9Eob�f� jFE�S��{�?�zZ���Bo�n�<7U����n)*J-S!Q