XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���V�FE�C��D�yG�g�8.3�{��ꒇ��Ud�To}�H���i]���2JZ7)����a
M�ηT�$I�1��`k��V�M�*4JzсzdF�#�z�<1�/��j�8ĵF�I����+h|�-ob3�>K��'@�g��s2�ٓ�*ͳ|Í2�.�K���k�w+�j*����f��]�se���m/�&�e��^��#؉.���Ɠ�R(���4�����	�~�u�jH����3�ZF/�ˇF�	@H�፼v����w�����wZ����˞*����QZl�*�*Q����~2y�C�4��Ҧ��m˺uN�C<�K�55C�+��R�.~��6�G7�M땠a�H�5@vH�?.���N<�=�b�S~D�^��WBwC/�f�m���q>Z�<=�մ�4Py��#ܝ )��NS�NU)U�M=/����K
H
��p���2��.���	�ޗ��Jj�d��0kq�+���}JWl���^����ΔmwHc�8�[���M�Ho,|�%�*h�$�ŒL�p���ԁp�&�e�ARڊJHY��sT�tR�;�kW �y8LO��-����gcu����M�d�l���me�:�|�W*p��]D�Y�X��B�]#�H��ݜȠzPH��%Q�z����L ��?����Ä*~W�f��j����Hlz�/f��<��������`��,EM=垟h���>��k&�Sc�\q��<��S�ͦϿ�"�R�� �T�XlxVHYEB    9efe    1be0�	��0�{�w�̡��E�}t�
�p���r�{��bS�`]Nf��T�`U��O�,����O�!��������TL唘i]��\�H:�=���ԝ�#<4�9-��j��ƀZ ��B�n��
(�#C~�H�,pq�ϣ
�]�MQE�$S_s{�)4_g�&y��<=�cr�ʍ\J梬-���CO�7��
��	kthD����4H��UC1q�b�ϥy$�-'��q[\A��:X�T]r���I\�
 `D�b�ߘb2��?�?����Ɠ��Z8�����	��Y�~oe�L��)sU�Ё{�\�����Vȳ�--�%!+��LN�Ϋ�|VN+��j�( �&ޖXw%u �lɑ����q�>��	����k��g���~�,J��p���!o��0��`K�=�a�8��=�����5���/�<F�,)�%_C5� /�ױ��58�}�e����+�23!3�D �#'��7���pB->�~o ➘<��^j�POT��X�����vު��dv�Ơ�o�x�������|��H��|f˾�1Չ�Yӫn�U��,C=��%I~9Ӿ]%*ԭ�H�埉dZW��w��d�����:�0`�=�/�@�o1�TŨ\~q�%�~(S�2�	F�s�=��E��xĬ=S�6�nJg�	���X��!�-�oS�Q ��#��rf�̢���F<7�����p����$���R`�/&�`_50G;?��P�[�ݝ���UQ��j�z�������4эU���.�x�z-�5�f;�1�jI�%�t|S4r��_�5�~m���6�>Fi�p��%�#C�}s��p����1T�K��'_O("����Y�3$��I���R��9��ND�J�3�՟���Yo�h�Z,�����6!��=.��#)C[{�2�O�B�(�泑�Ֆ~���+D�\ǩ�/Hk�0�V���M�>F��]�g��j5�
U��A b�#-y��V{.H
�RB���+�D��2v�"���`�Tn�@�����Ha��P�0Wa����3�ץ'͝�u��,X�{���^�p�ac����9/�����y<�q�C�Td�2LE�j��|�b;����8`r�%UC�O�שJ0�O�<[��J:5�����X�L�ǆ4? 2����bd��6�QO?�U��}1���7�]������փ~W�H�g��Ity�5\i2;;DQC2Kނ~υCw�f̉�l��zΒ�0��¿/�B{��8G��"�&*��.��<[������$?�6�MJ�3����E}zU�	����\�H7Ȏ�����:4q9��{�ǃ����ւVG[܁&ۡ5���9'`k�Z��S���؞�r6� 9L� 3�f�%���@D>� e�{[�H�)p��5G��PVh]���/P_��=C�aY���o��]e��H��C^Dc�n���z4C�DJ�y�Q�(o3PSu��d�Hf�r6 ��c�!Dv,0=�s�.~���]��A�ǬXNc睖ԇ~�����1��ND`���t��F�e��?�����:�Ԗ�O�ךN��;����D�~J�Ð�@[A8gG%��!�a���?R1MעJ^>� ��TJ愉)h����]���������E��^�&��W�І����o�}w�Y���]͝!����h�l�{�
å���vY��  [V'�ZS�����|����:�~�`��j<3'u{�:�~(Pd��x���l��ܬi4��|!,�r�W�wc���/��=Gjм�͚�f�W��[D��4��0�+�:��|^�*���d��%�C����џ�ք))���i�K}tˠVY���ë�G|n8ʚ��h�[��W�m?����u�!����5�`�>~��?��t�lA��:��?!s���oO�)O�0�uBAePK'���f:���72��&�ѽ��yI�:��	,�8W�b��i|��Q��q���b؞�j� w�
?�]C��$ŋ\m��OU]�}C��n�E�geJ�OôO/��<���Z�&�C��f���Eˣ���OD�E3���W�cSBȼ�����0��n�e󕧏�u�f���>�h������CE�Sڿ_$U��	Q(�ռ����M�k��=]�v�5��H';�]8xM�?��j򊓐�1:�@dNr��D��m�5S�)��>߫�Г�۝�����S�i�\v ���[��V���1b��?����2��=���R�ţ ZN_������\�r�A��������}urҬL�^���T5�˭�X��$���ğ	5Z��B�GD��R�X����:|����j����C#�(kcmr�n1-����Ց
>�WT��@�v��������A��W{�.�����k�nNǀ<cw$�\ie�"�z6Y��%o&�Kں�����̃��PyiGkC�����Α�5���y�!2�L�H(k 	$)�u��ֵ��@���Y��g�g�:���F��F��6�	�.(p��z�C}��7�Ɏ�C=�B���Г&*�~��^7f��ɒ+�K����n��L�b����H�x۳�CG�"�1u�\����#�Y��̋+Ѣ�թ�4U� ��B���"i� y�X����\���[�N}���#�z� ��~d9r�ƹ%��Q҉����%����oV_}�x��.�ͅay!�����v��$T(6�,��{	� �H�<�Z��)�n �ײ,f�
�ϰ�&�;ۨ�,���X�X�H�Ona4?�S������+��1^�c�,�i���?"R�Yi���<�sKO�j�����ܘ�Y;,��
uQ�qp��$���Uؕ&��9߳+��i�`�-A���\�-�
�0�Ͷ����J��산�;Z�������i�t����'�������i{��YQ)�p�L� �1Ri�,�y"�[k$H�Ė��')C[0K;ە�}����E$%�)<h��}���Q>՚U�H٩�"� �6�����������4d� �ѩѱЈ�wr�빪��R���G؏�t�kУ��b�_�N�.�dP1e2��	�ZHz�<S�@�.�����5��l����1�3�/��`g��������Wȳ<�"��aa$�`꾾���,�O� W��@����"$����v�d��t������Ζ� �9Frs�����h	���A֡F�虢�c�Մp��Z���BB<p�:vqE(?r�oԓm`ս|9Ux ۴�������� �䐗���7U(�&5�V����/� V�[x��ŠX��uu�$�=MdV�Jh�V	ӛ����WB�=|�K]��0Lˢ���ԑ	���3�4�����"@0aH�u˴�.`D|#�S ��� �?3�#WƮ�����R;��u�1 � y�oO(kK�fЋj��Қo�EuYLHA��kl��M�hJ�������?���b�L9!��_tY� � Zu�Ɍ�(+��Q��
[�K�J����a����(�qiZ�n!:��h��,�FA��!��a���鍜���x,�#�E��m6��ؒ7�K�Z���_؇�-Y�غwٔ�W�e�b�s�Yi��U'^�������ֈ��*����.�7io�(���[Z�h�6���$f�
�]�ƅ�n�S��F�M���J��$�5�:w!`O��"���~�����pp�y����h�eJ_���@�����G��lV	?F���C�FG`(��K:��5��ǅd�!vP�@n!~�y� ��T�/��ű���ۯ������2�+��8D���w�0_��}|6,���KB���%�J�p�lC��$�o��&g��hL�k����QoX0��,�AR��~h;bW�~�"��mH~���OzWO�쮓�r�6P<Q�l��׾�Pa��;E��Xa|�/[�q���V�-l���ʢ[�x徟5~��Q�/�m���ݭ�6a 	KRؒp4K}I\Z&
vW�-�4��ʇ�6�]�p�����!�h/�jW�yR������x�{����@q�,�o�L�v/V�{�w��w�����t�t����LK�������E��9�!ׂ�/\���I'��.N�L�
�]Lȟ����Z�"�CS��=�!���zp�TW�7�4���Gr�Nvw C��N�I�@���C��	�Dj��t6iD��0\��\2*@R�9���3�E;�9r��3 �D��J'�">�9xe�X�Zר���!d_����+x0����Z�O�:�^J��s��HԪ��H����t�F��Eؒ�Ӯ蛾lZ��D!%r~W�#�jZ��V93t�����{k��&M�=���edD���X|�J��(7)@ˮ������`��b�\�D�
��n_�%�q��G�إ�dN(o҈���#�,�B>Sq��>>��]�ҮE�]���R�#b�lZ�G�4?����"ƨ��cߜ����t��%%6V:2yf!}Eo4|�x'ŜuEd�oDqQ�eo@�	���*V��-g��8u����K�gҦj[!�ės�0n*����8DL3W�D�	0:Jl��a
���eL�����,Nx7���9�� }�{z��� b!i����Y"�L�a��j͈�"L���|,�Z�Ea�sL�K7t��9��+�~���b�1瞎B���VC�������i�g���;+c���?Bb[�|)��mwrKT��Ik��C �����J��<��U���Ocӈb��u�<S�@u����c��"�7p6<g�J��� `y�h{Qб�>�h��D�0�R�'&��I��Z�_=��H � A�������1�{�o���R|��� �����#�1���y�����!�ƶ��#7����>o��cat�}�+s��9	r���*l��8a^�7v;f5��ԅ� n3���;�5(�OH��D��K1��Q�3b�!�5e
�+�&�E/d�J<�1(1�N��سDТQ�z��#'��R����I��C�dȦ]��x�4��u�,$s�R�^K9amo܈J�
�#��$O?]�=p��T��k ��u�3�Ĩ��b~�|y��c}���傎���-ު(���u�L���q3�r��6IO��I�+R�r��T����Uڒ����=+˽�g��d��ܢ���W�����z��~y����G#� rn�;�O�����u�����%@�40� �����pO�=�,�f��B9�AUY��v�8s�׆O�y�ܶG�1�E����FJGk�m� p��1����3�x�$&�vw�d��O�L/�{;'���¢E����?ق��D���Mi ��\e�=�A��pr��veR�Y�9%�s�I@�IT��ͪ(i@�ҏ��F	�X,�n�~�T���'��6Olk��yu���6��
Z����B6t����\/3��ڶ��Z�^W��g�w�+�B��3�8 5 �s�4� ��:c���.k&\3<��0�������N|����@��:[��*��&Yj0��W)"̺,�a���wH�'~�u�AY�	XOד�|n��r��з�|�����{�@��~�sm+q�W�3Z���51^gS�=�b�c7���~B�Z��<�!E��X�j��맇�#G�k`x�X@� ,��
�C#�q�R�>lACg%NW�0��SPo�������r�J+����!F �[9nރ*W����+�q�ʀh��Q� -ՄQ.��Bi�e��a�z ��"�'D��W�K�q��e7՗}�|@���M���(qs|p*�,���@1@���;AhNA��I�}��c���2U�*P�bAP cu�5A�κ�n�r�GimC��ث>���$Rg�7�W�^����{�WQG(������$���U�<V�7A���攞	�,R-�_������0�;�k��l�%W7Jţϳ=��lz����b�г���ЧG�{+ҳ\8�e��Y�vW�n�@���0�=ޒ���Gn[�&M�?z�iCZ��I.K8|��:�#���\������f@���8���Jf?$���W<W�e#؂'���Vs�-�\`�>%���5������S��j.sx�O'�����Wg*-�O�3=�b�ّ�p��(�<o^mȓ<�PAt��
	av8J��L&���Z�n�s��:�IK�k{[q�H���$\m���XՒ��h��0(���s�`: 	���/���
"��E��sa.�F������!R'�p^-ݴ�kXm0��$)s/³\Q�W���e>��h����ڂ� ���'#�&B-M�~ya�(�2���v�v�4-���vf�kʄ����Wn��F@��:�sq���ƴ����-E������]��g|J��"��T1�{&�DNǛ���^S�U& ʁ@q<;̿ �|��+SR<������Vh5l'��C�$�Ͱ�kD�+$U_4S����)�{��y5��+��#�/��Yr��{�lܶ4���
�;�!�U��X��	��aB�2�����\�d�r䝧�����d�����3�[7_��xMy�l�(�h�/�7V0��L]Z�\��9 ~�N�E����s�IE��ʇ�y�R�N�FW�F��wmS1:f{�ɧ��>����Uq��$�az{ż�]x�I��s�Q�!Lk>rh}���{�듊W�9S�`q��\�ࡗl�d��q�`oA'��֪'%�um%�+Dcy��q�P�����ߑ^Q<�n�B�gd��x��9!�{
��*ce}6@���9֤���RW<�vM���+@�Ζ��m�*��\=ƾj�_�I�$�Jjo������Y��S��i�>��Q�sؼg���9偑�@{���$k	��JB����ϛ^'�"G�&���߂p!lVeB��Q6a�gq4G�ae��b)�7��j�odl��t b�%���g��D��u�o���ܪtL�4T�X!
�#�G�"{o��Qդ�B>���d_������Q7��}�9��}�����턮��BK���B��?�q�a-�"�M0���,A1�e��\�e��P�A\%f@��pm̉�